module CRat(
  input        clock,
               reset,
  input  [4:0] io_rj_0,
               io_rj_1,
               io_rj_2,
               io_rj_3,
               io_rk_0,
               io_rk_1,
               io_rk_2,
               io_rk_3,
               io_rd_0,
               io_rd_1,
               io_rd_2,
               io_rd_3,
  input        io_rd_valid_0,
               io_rd_valid_1,
               io_rd_valid_2,
               io_rd_valid_3,
  input  [5:0] io_alloc_preg_0,
               io_alloc_preg_1,
               io_alloc_preg_2,
               io_alloc_preg_3,
  input        io_arch_rat_0,
               io_arch_rat_1,
               io_arch_rat_2,
               io_arch_rat_3,
               io_arch_rat_4,
               io_arch_rat_5,
               io_arch_rat_6,
               io_arch_rat_7,
               io_arch_rat_8,
               io_arch_rat_9,
               io_arch_rat_10,
               io_arch_rat_11,
               io_arch_rat_12,
               io_arch_rat_13,
               io_arch_rat_14,
               io_arch_rat_15,
               io_arch_rat_16,
               io_arch_rat_17,
               io_arch_rat_18,
               io_arch_rat_19,
               io_arch_rat_20,
               io_arch_rat_21,
               io_arch_rat_22,
               io_arch_rat_23,
               io_arch_rat_24,
               io_arch_rat_25,
               io_arch_rat_26,
               io_arch_rat_27,
               io_arch_rat_28,
               io_arch_rat_29,
               io_arch_rat_30,
               io_arch_rat_31,
               io_arch_rat_32,
               io_arch_rat_33,
               io_arch_rat_34,
               io_arch_rat_35,
               io_arch_rat_36,
               io_arch_rat_37,
               io_arch_rat_38,
               io_arch_rat_39,
               io_arch_rat_40,
               io_arch_rat_41,
               io_arch_rat_42,
               io_arch_rat_43,
               io_arch_rat_44,
               io_arch_rat_45,
               io_arch_rat_46,
               io_arch_rat_47,
               io_arch_rat_48,
               io_arch_rat_49,
               io_arch_rat_50,
               io_arch_rat_51,
               io_arch_rat_52,
               io_arch_rat_53,
               io_arch_rat_54,
               io_arch_rat_55,
               io_arch_rat_56,
               io_arch_rat_57,
               io_arch_rat_58,
               io_arch_rat_59,
               io_arch_rat_60,
               io_arch_rat_61,
               io_arch_rat_62,
               io_arch_rat_63,
               io_predict_fail,
  output [5:0] io_prj_0,
               io_prj_1,
               io_prj_2,
               io_prj_3,
               io_prk_0,
               io_prk_1,
               io_prk_2,
               io_prk_3,
               io_pprd_0,
               io_pprd_1,
               io_pprd_2,
               io_pprd_3
);

  reg         crat_0_valid;
  reg  [4:0]  crat_0_lr;
  reg         crat_1_valid;
  reg  [4:0]  crat_1_lr;
  reg         crat_2_valid;
  reg  [4:0]  crat_2_lr;
  reg         crat_3_valid;
  reg  [4:0]  crat_3_lr;
  reg         crat_4_valid;
  reg  [4:0]  crat_4_lr;
  reg         crat_5_valid;
  reg  [4:0]  crat_5_lr;
  reg         crat_6_valid;
  reg  [4:0]  crat_6_lr;
  reg         crat_7_valid;
  reg  [4:0]  crat_7_lr;
  reg         crat_8_valid;
  reg  [4:0]  crat_8_lr;
  reg         crat_9_valid;
  reg  [4:0]  crat_9_lr;
  reg         crat_10_valid;
  reg  [4:0]  crat_10_lr;
  reg         crat_11_valid;
  reg  [4:0]  crat_11_lr;
  reg         crat_12_valid;
  reg  [4:0]  crat_12_lr;
  reg         crat_13_valid;
  reg  [4:0]  crat_13_lr;
  reg         crat_14_valid;
  reg  [4:0]  crat_14_lr;
  reg         crat_15_valid;
  reg  [4:0]  crat_15_lr;
  reg         crat_16_valid;
  reg  [4:0]  crat_16_lr;
  reg         crat_17_valid;
  reg  [4:0]  crat_17_lr;
  reg         crat_18_valid;
  reg  [4:0]  crat_18_lr;
  reg         crat_19_valid;
  reg  [4:0]  crat_19_lr;
  reg         crat_20_valid;
  reg  [4:0]  crat_20_lr;
  reg         crat_21_valid;
  reg  [4:0]  crat_21_lr;
  reg         crat_22_valid;
  reg  [4:0]  crat_22_lr;
  reg         crat_23_valid;
  reg  [4:0]  crat_23_lr;
  reg         crat_24_valid;
  reg  [4:0]  crat_24_lr;
  reg         crat_25_valid;
  reg  [4:0]  crat_25_lr;
  reg         crat_26_valid;
  reg  [4:0]  crat_26_lr;
  reg         crat_27_valid;
  reg  [4:0]  crat_27_lr;
  reg         crat_28_valid;
  reg  [4:0]  crat_28_lr;
  reg         crat_29_valid;
  reg  [4:0]  crat_29_lr;
  reg         crat_30_valid;
  reg  [4:0]  crat_30_lr;
  reg         crat_31_valid;
  reg  [4:0]  crat_31_lr;
  reg         crat_32_valid;
  reg  [4:0]  crat_32_lr;
  reg         crat_33_valid;
  reg  [4:0]  crat_33_lr;
  reg         crat_34_valid;
  reg  [4:0]  crat_34_lr;
  reg         crat_35_valid;
  reg  [4:0]  crat_35_lr;
  reg         crat_36_valid;
  reg  [4:0]  crat_36_lr;
  reg         crat_37_valid;
  reg  [4:0]  crat_37_lr;
  reg         crat_38_valid;
  reg  [4:0]  crat_38_lr;
  reg         crat_39_valid;
  reg  [4:0]  crat_39_lr;
  reg         crat_40_valid;
  reg  [4:0]  crat_40_lr;
  reg         crat_41_valid;
  reg  [4:0]  crat_41_lr;
  reg         crat_42_valid;
  reg  [4:0]  crat_42_lr;
  reg         crat_43_valid;
  reg  [4:0]  crat_43_lr;
  reg         crat_44_valid;
  reg  [4:0]  crat_44_lr;
  reg         crat_45_valid;
  reg  [4:0]  crat_45_lr;
  reg         crat_46_valid;
  reg  [4:0]  crat_46_lr;
  reg         crat_47_valid;
  reg  [4:0]  crat_47_lr;
  reg         crat_48_valid;
  reg  [4:0]  crat_48_lr;
  reg         crat_49_valid;
  reg  [4:0]  crat_49_lr;
  reg         crat_50_valid;
  reg  [4:0]  crat_50_lr;
  reg         crat_51_valid;
  reg  [4:0]  crat_51_lr;
  reg         crat_52_valid;
  reg  [4:0]  crat_52_lr;
  reg         crat_53_valid;
  reg  [4:0]  crat_53_lr;
  reg         crat_54_valid;
  reg  [4:0]  crat_54_lr;
  reg         crat_55_valid;
  reg  [4:0]  crat_55_lr;
  reg         crat_56_valid;
  reg  [4:0]  crat_56_lr;
  reg         crat_57_valid;
  reg  [4:0]  crat_57_lr;
  reg         crat_58_valid;
  reg  [4:0]  crat_58_lr;
  reg         crat_59_valid;
  reg  [4:0]  crat_59_lr;
  reg         crat_60_valid;
  reg  [4:0]  crat_60_lr;
  reg         crat_61_valid;
  reg  [4:0]  crat_61_lr;
  reg         crat_62_valid;
  reg  [4:0]  crat_62_lr;
  reg         crat_63_valid;
  reg  [4:0]  crat_63_lr;
  wire        rj_hit_oh_0_33 = crat_33_valid & crat_33_lr == io_rj_0;
  wire        rk_hit_oh_0_33 = crat_33_valid & crat_33_lr == io_rk_0;
  wire        rd_hit_oh_0_33 = crat_33_valid & crat_33_lr == io_rd_0;
  wire        rj_hit_oh_0_34 = crat_34_valid & crat_34_lr == io_rj_0;
  wire        rk_hit_oh_0_34 = crat_34_valid & crat_34_lr == io_rk_0;
  wire        rd_hit_oh_0_34 = crat_34_valid & crat_34_lr == io_rd_0;
  wire        rj_hit_oh_0_35 = crat_35_valid & crat_35_lr == io_rj_0;
  wire        rk_hit_oh_0_35 = crat_35_valid & crat_35_lr == io_rk_0;
  wire        rd_hit_oh_0_35 = crat_35_valid & crat_35_lr == io_rd_0;
  wire        rj_hit_oh_0_36 = crat_36_valid & crat_36_lr == io_rj_0;
  wire        rk_hit_oh_0_36 = crat_36_valid & crat_36_lr == io_rk_0;
  wire        rd_hit_oh_0_36 = crat_36_valid & crat_36_lr == io_rd_0;
  wire        rj_hit_oh_0_37 = crat_37_valid & crat_37_lr == io_rj_0;
  wire        rk_hit_oh_0_37 = crat_37_valid & crat_37_lr == io_rk_0;
  wire        rd_hit_oh_0_37 = crat_37_valid & crat_37_lr == io_rd_0;
  wire        rj_hit_oh_0_38 = crat_38_valid & crat_38_lr == io_rj_0;
  wire        rk_hit_oh_0_38 = crat_38_valid & crat_38_lr == io_rk_0;
  wire        rd_hit_oh_0_38 = crat_38_valid & crat_38_lr == io_rd_0;
  wire        rj_hit_oh_0_39 = crat_39_valid & crat_39_lr == io_rj_0;
  wire        rk_hit_oh_0_39 = crat_39_valid & crat_39_lr == io_rk_0;
  wire        rd_hit_oh_0_39 = crat_39_valid & crat_39_lr == io_rd_0;
  wire        rj_hit_oh_0_40 = crat_40_valid & crat_40_lr == io_rj_0;
  wire        rk_hit_oh_0_40 = crat_40_valid & crat_40_lr == io_rk_0;
  wire        rd_hit_oh_0_40 = crat_40_valid & crat_40_lr == io_rd_0;
  wire        rj_hit_oh_0_41 = crat_41_valid & crat_41_lr == io_rj_0;
  wire        rk_hit_oh_0_41 = crat_41_valid & crat_41_lr == io_rk_0;
  wire        rd_hit_oh_0_41 = crat_41_valid & crat_41_lr == io_rd_0;
  wire        rj_hit_oh_0_42 = crat_42_valid & crat_42_lr == io_rj_0;
  wire        rk_hit_oh_0_42 = crat_42_valid & crat_42_lr == io_rk_0;
  wire        rd_hit_oh_0_42 = crat_42_valid & crat_42_lr == io_rd_0;
  wire        rj_hit_oh_0_43 = crat_43_valid & crat_43_lr == io_rj_0;
  wire        rk_hit_oh_0_43 = crat_43_valid & crat_43_lr == io_rk_0;
  wire        rd_hit_oh_0_43 = crat_43_valid & crat_43_lr == io_rd_0;
  wire        rj_hit_oh_0_44 = crat_44_valid & crat_44_lr == io_rj_0;
  wire        rk_hit_oh_0_44 = crat_44_valid & crat_44_lr == io_rk_0;
  wire        rd_hit_oh_0_44 = crat_44_valid & crat_44_lr == io_rd_0;
  wire        rj_hit_oh_0_45 = crat_45_valid & crat_45_lr == io_rj_0;
  wire        rk_hit_oh_0_45 = crat_45_valid & crat_45_lr == io_rk_0;
  wire        rd_hit_oh_0_45 = crat_45_valid & crat_45_lr == io_rd_0;
  wire        rj_hit_oh_0_46 = crat_46_valid & crat_46_lr == io_rj_0;
  wire        rk_hit_oh_0_46 = crat_46_valid & crat_46_lr == io_rk_0;
  wire        rd_hit_oh_0_46 = crat_46_valid & crat_46_lr == io_rd_0;
  wire        rj_hit_oh_0_47 = crat_47_valid & crat_47_lr == io_rj_0;
  wire        rk_hit_oh_0_47 = crat_47_valid & crat_47_lr == io_rk_0;
  wire        rd_hit_oh_0_47 = crat_47_valid & crat_47_lr == io_rd_0;
  wire        rj_hit_oh_0_48 = crat_48_valid & crat_48_lr == io_rj_0;
  wire        rk_hit_oh_0_48 = crat_48_valid & crat_48_lr == io_rk_0;
  wire        rd_hit_oh_0_48 = crat_48_valid & crat_48_lr == io_rd_0;
  wire        rj_hit_oh_0_49 = crat_49_valid & crat_49_lr == io_rj_0;
  wire        rk_hit_oh_0_49 = crat_49_valid & crat_49_lr == io_rk_0;
  wire        rd_hit_oh_0_49 = crat_49_valid & crat_49_lr == io_rd_0;
  wire        rj_hit_oh_0_50 = crat_50_valid & crat_50_lr == io_rj_0;
  wire        rk_hit_oh_0_50 = crat_50_valid & crat_50_lr == io_rk_0;
  wire        rd_hit_oh_0_50 = crat_50_valid & crat_50_lr == io_rd_0;
  wire        rj_hit_oh_0_51 = crat_51_valid & crat_51_lr == io_rj_0;
  wire        rk_hit_oh_0_51 = crat_51_valid & crat_51_lr == io_rk_0;
  wire        rd_hit_oh_0_51 = crat_51_valid & crat_51_lr == io_rd_0;
  wire        rj_hit_oh_0_52 = crat_52_valid & crat_52_lr == io_rj_0;
  wire        rk_hit_oh_0_52 = crat_52_valid & crat_52_lr == io_rk_0;
  wire        rd_hit_oh_0_52 = crat_52_valid & crat_52_lr == io_rd_0;
  wire        rj_hit_oh_0_53 = crat_53_valid & crat_53_lr == io_rj_0;
  wire        rk_hit_oh_0_53 = crat_53_valid & crat_53_lr == io_rk_0;
  wire        rd_hit_oh_0_53 = crat_53_valid & crat_53_lr == io_rd_0;
  wire        rj_hit_oh_0_54 = crat_54_valid & crat_54_lr == io_rj_0;
  wire        rk_hit_oh_0_54 = crat_54_valid & crat_54_lr == io_rk_0;
  wire        rd_hit_oh_0_54 = crat_54_valid & crat_54_lr == io_rd_0;
  wire        rj_hit_oh_0_55 = crat_55_valid & crat_55_lr == io_rj_0;
  wire        rk_hit_oh_0_55 = crat_55_valid & crat_55_lr == io_rk_0;
  wire        rd_hit_oh_0_55 = crat_55_valid & crat_55_lr == io_rd_0;
  wire        rj_hit_oh_0_56 = crat_56_valid & crat_56_lr == io_rj_0;
  wire        rk_hit_oh_0_56 = crat_56_valid & crat_56_lr == io_rk_0;
  wire        rd_hit_oh_0_56 = crat_56_valid & crat_56_lr == io_rd_0;
  wire        rj_hit_oh_0_57 = crat_57_valid & crat_57_lr == io_rj_0;
  wire        rk_hit_oh_0_57 = crat_57_valid & crat_57_lr == io_rk_0;
  wire        rd_hit_oh_0_57 = crat_57_valid & crat_57_lr == io_rd_0;
  wire        rj_hit_oh_0_58 = crat_58_valid & crat_58_lr == io_rj_0;
  wire        rk_hit_oh_0_58 = crat_58_valid & crat_58_lr == io_rk_0;
  wire        rd_hit_oh_0_58 = crat_58_valid & crat_58_lr == io_rd_0;
  wire        rj_hit_oh_0_59 = crat_59_valid & crat_59_lr == io_rj_0;
  wire        rk_hit_oh_0_59 = crat_59_valid & crat_59_lr == io_rk_0;
  wire        rd_hit_oh_0_59 = crat_59_valid & crat_59_lr == io_rd_0;
  wire        rj_hit_oh_0_60 = crat_60_valid & crat_60_lr == io_rj_0;
  wire        rk_hit_oh_0_60 = crat_60_valid & crat_60_lr == io_rk_0;
  wire        rd_hit_oh_0_60 = crat_60_valid & crat_60_lr == io_rd_0;
  wire        rj_hit_oh_0_61 = crat_61_valid & crat_61_lr == io_rj_0;
  wire        rk_hit_oh_0_61 = crat_61_valid & crat_61_lr == io_rk_0;
  wire        rd_hit_oh_0_61 = crat_61_valid & crat_61_lr == io_rd_0;
  wire        rj_hit_oh_0_62 = crat_62_valid & crat_62_lr == io_rj_0;
  wire        rk_hit_oh_0_62 = crat_62_valid & crat_62_lr == io_rk_0;
  wire        rd_hit_oh_0_62 = crat_62_valid & crat_62_lr == io_rd_0;
  wire        rj_hit_oh_0_63 = crat_63_valid & crat_63_lr == io_rj_0;
  wire        rk_hit_oh_0_63 = crat_63_valid & crat_63_lr == io_rk_0;
  wire        rd_hit_oh_0_63 = crat_63_valid & crat_63_lr == io_rd_0;
  wire [30:0] _io_prj_0_T_1073 =
    {rj_hit_oh_0_63,
     rj_hit_oh_0_62,
     rj_hit_oh_0_61,
     rj_hit_oh_0_60,
     rj_hit_oh_0_59,
     rj_hit_oh_0_58,
     rj_hit_oh_0_57,
     rj_hit_oh_0_56,
     rj_hit_oh_0_55,
     rj_hit_oh_0_54,
     rj_hit_oh_0_53,
     rj_hit_oh_0_52,
     rj_hit_oh_0_51,
     rj_hit_oh_0_50,
     rj_hit_oh_0_49,
     rj_hit_oh_0_48,
     rj_hit_oh_0_47,
     rj_hit_oh_0_46,
     rj_hit_oh_0_45,
     rj_hit_oh_0_44,
     rj_hit_oh_0_43,
     rj_hit_oh_0_42,
     rj_hit_oh_0_41,
     rj_hit_oh_0_40,
     rj_hit_oh_0_39,
     rj_hit_oh_0_38,
     rj_hit_oh_0_37,
     rj_hit_oh_0_36,
     rj_hit_oh_0_35,
     rj_hit_oh_0_34,
     rj_hit_oh_0_33}
    | {crat_31_valid & crat_31_lr == io_rj_0,
       crat_30_valid & crat_30_lr == io_rj_0,
       crat_29_valid & crat_29_lr == io_rj_0,
       crat_28_valid & crat_28_lr == io_rj_0,
       crat_27_valid & crat_27_lr == io_rj_0,
       crat_26_valid & crat_26_lr == io_rj_0,
       crat_25_valid & crat_25_lr == io_rj_0,
       crat_24_valid & crat_24_lr == io_rj_0,
       crat_23_valid & crat_23_lr == io_rj_0,
       crat_22_valid & crat_22_lr == io_rj_0,
       crat_21_valid & crat_21_lr == io_rj_0,
       crat_20_valid & crat_20_lr == io_rj_0,
       crat_19_valid & crat_19_lr == io_rj_0,
       crat_18_valid & crat_18_lr == io_rj_0,
       crat_17_valid & crat_17_lr == io_rj_0,
       crat_16_valid & crat_16_lr == io_rj_0,
       crat_15_valid & crat_15_lr == io_rj_0,
       crat_14_valid & crat_14_lr == io_rj_0,
       crat_13_valid & crat_13_lr == io_rj_0,
       crat_12_valid & crat_12_lr == io_rj_0,
       crat_11_valid & crat_11_lr == io_rj_0,
       crat_10_valid & crat_10_lr == io_rj_0,
       crat_9_valid & crat_9_lr == io_rj_0,
       crat_8_valid & crat_8_lr == io_rj_0,
       crat_7_valid & crat_7_lr == io_rj_0,
       crat_6_valid & crat_6_lr == io_rj_0,
       crat_5_valid & crat_5_lr == io_rj_0,
       crat_4_valid & crat_4_lr == io_rj_0,
       crat_3_valid & crat_3_lr == io_rj_0,
       crat_2_valid & crat_2_lr == io_rj_0,
       crat_1_valid & crat_1_lr == io_rj_0};
  wire [14:0] _io_prj_0_T_1075 = _io_prj_0_T_1073[30:16] | _io_prj_0_T_1073[14:0];
  wire [6:0]  _io_prj_0_T_1077 = _io_prj_0_T_1075[14:8] | _io_prj_0_T_1075[6:0];
  wire [2:0]  _io_prj_0_T_1079 = _io_prj_0_T_1077[6:4] | _io_prj_0_T_1077[2:0];
  wire [30:0] _io_prk_0_T_1073 =
    {rk_hit_oh_0_63,
     rk_hit_oh_0_62,
     rk_hit_oh_0_61,
     rk_hit_oh_0_60,
     rk_hit_oh_0_59,
     rk_hit_oh_0_58,
     rk_hit_oh_0_57,
     rk_hit_oh_0_56,
     rk_hit_oh_0_55,
     rk_hit_oh_0_54,
     rk_hit_oh_0_53,
     rk_hit_oh_0_52,
     rk_hit_oh_0_51,
     rk_hit_oh_0_50,
     rk_hit_oh_0_49,
     rk_hit_oh_0_48,
     rk_hit_oh_0_47,
     rk_hit_oh_0_46,
     rk_hit_oh_0_45,
     rk_hit_oh_0_44,
     rk_hit_oh_0_43,
     rk_hit_oh_0_42,
     rk_hit_oh_0_41,
     rk_hit_oh_0_40,
     rk_hit_oh_0_39,
     rk_hit_oh_0_38,
     rk_hit_oh_0_37,
     rk_hit_oh_0_36,
     rk_hit_oh_0_35,
     rk_hit_oh_0_34,
     rk_hit_oh_0_33}
    | {crat_31_valid & crat_31_lr == io_rk_0,
       crat_30_valid & crat_30_lr == io_rk_0,
       crat_29_valid & crat_29_lr == io_rk_0,
       crat_28_valid & crat_28_lr == io_rk_0,
       crat_27_valid & crat_27_lr == io_rk_0,
       crat_26_valid & crat_26_lr == io_rk_0,
       crat_25_valid & crat_25_lr == io_rk_0,
       crat_24_valid & crat_24_lr == io_rk_0,
       crat_23_valid & crat_23_lr == io_rk_0,
       crat_22_valid & crat_22_lr == io_rk_0,
       crat_21_valid & crat_21_lr == io_rk_0,
       crat_20_valid & crat_20_lr == io_rk_0,
       crat_19_valid & crat_19_lr == io_rk_0,
       crat_18_valid & crat_18_lr == io_rk_0,
       crat_17_valid & crat_17_lr == io_rk_0,
       crat_16_valid & crat_16_lr == io_rk_0,
       crat_15_valid & crat_15_lr == io_rk_0,
       crat_14_valid & crat_14_lr == io_rk_0,
       crat_13_valid & crat_13_lr == io_rk_0,
       crat_12_valid & crat_12_lr == io_rk_0,
       crat_11_valid & crat_11_lr == io_rk_0,
       crat_10_valid & crat_10_lr == io_rk_0,
       crat_9_valid & crat_9_lr == io_rk_0,
       crat_8_valid & crat_8_lr == io_rk_0,
       crat_7_valid & crat_7_lr == io_rk_0,
       crat_6_valid & crat_6_lr == io_rk_0,
       crat_5_valid & crat_5_lr == io_rk_0,
       crat_4_valid & crat_4_lr == io_rk_0,
       crat_3_valid & crat_3_lr == io_rk_0,
       crat_2_valid & crat_2_lr == io_rk_0,
       crat_1_valid & crat_1_lr == io_rk_0};
  wire [14:0] _io_prk_0_T_1075 = _io_prk_0_T_1073[30:16] | _io_prk_0_T_1073[14:0];
  wire [6:0]  _io_prk_0_T_1077 = _io_prk_0_T_1075[14:8] | _io_prk_0_T_1075[6:0];
  wire [2:0]  _io_prk_0_T_1079 = _io_prk_0_T_1077[6:4] | _io_prk_0_T_1077[2:0];
  wire [30:0] _io_pprd_0_T_1073 =
    {rd_hit_oh_0_63,
     rd_hit_oh_0_62,
     rd_hit_oh_0_61,
     rd_hit_oh_0_60,
     rd_hit_oh_0_59,
     rd_hit_oh_0_58,
     rd_hit_oh_0_57,
     rd_hit_oh_0_56,
     rd_hit_oh_0_55,
     rd_hit_oh_0_54,
     rd_hit_oh_0_53,
     rd_hit_oh_0_52,
     rd_hit_oh_0_51,
     rd_hit_oh_0_50,
     rd_hit_oh_0_49,
     rd_hit_oh_0_48,
     rd_hit_oh_0_47,
     rd_hit_oh_0_46,
     rd_hit_oh_0_45,
     rd_hit_oh_0_44,
     rd_hit_oh_0_43,
     rd_hit_oh_0_42,
     rd_hit_oh_0_41,
     rd_hit_oh_0_40,
     rd_hit_oh_0_39,
     rd_hit_oh_0_38,
     rd_hit_oh_0_37,
     rd_hit_oh_0_36,
     rd_hit_oh_0_35,
     rd_hit_oh_0_34,
     rd_hit_oh_0_33}
    | {crat_31_valid & crat_31_lr == io_rd_0,
       crat_30_valid & crat_30_lr == io_rd_0,
       crat_29_valid & crat_29_lr == io_rd_0,
       crat_28_valid & crat_28_lr == io_rd_0,
       crat_27_valid & crat_27_lr == io_rd_0,
       crat_26_valid & crat_26_lr == io_rd_0,
       crat_25_valid & crat_25_lr == io_rd_0,
       crat_24_valid & crat_24_lr == io_rd_0,
       crat_23_valid & crat_23_lr == io_rd_0,
       crat_22_valid & crat_22_lr == io_rd_0,
       crat_21_valid & crat_21_lr == io_rd_0,
       crat_20_valid & crat_20_lr == io_rd_0,
       crat_19_valid & crat_19_lr == io_rd_0,
       crat_18_valid & crat_18_lr == io_rd_0,
       crat_17_valid & crat_17_lr == io_rd_0,
       crat_16_valid & crat_16_lr == io_rd_0,
       crat_15_valid & crat_15_lr == io_rd_0,
       crat_14_valid & crat_14_lr == io_rd_0,
       crat_13_valid & crat_13_lr == io_rd_0,
       crat_12_valid & crat_12_lr == io_rd_0,
       crat_11_valid & crat_11_lr == io_rd_0,
       crat_10_valid & crat_10_lr == io_rd_0,
       crat_9_valid & crat_9_lr == io_rd_0,
       crat_8_valid & crat_8_lr == io_rd_0,
       crat_7_valid & crat_7_lr == io_rd_0,
       crat_6_valid & crat_6_lr == io_rd_0,
       crat_5_valid & crat_5_lr == io_rd_0,
       crat_4_valid & crat_4_lr == io_rd_0,
       crat_3_valid & crat_3_lr == io_rd_0,
       crat_2_valid & crat_2_lr == io_rd_0,
       crat_1_valid & crat_1_lr == io_rd_0};
  wire [14:0] _io_pprd_0_T_1075 = _io_pprd_0_T_1073[30:16] | _io_pprd_0_T_1073[14:0];
  wire [6:0]  _io_pprd_0_T_1077 = _io_pprd_0_T_1075[14:8] | _io_pprd_0_T_1075[6:0];
  wire [2:0]  _io_pprd_0_T_1079 = _io_pprd_0_T_1077[6:4] | _io_pprd_0_T_1077[2:0];
  wire [5:0]  _io_pprd_0_output =
    {|{rd_hit_oh_0_63,
       rd_hit_oh_0_62,
       rd_hit_oh_0_61,
       rd_hit_oh_0_60,
       rd_hit_oh_0_59,
       rd_hit_oh_0_58,
       rd_hit_oh_0_57,
       rd_hit_oh_0_56,
       rd_hit_oh_0_55,
       rd_hit_oh_0_54,
       rd_hit_oh_0_53,
       rd_hit_oh_0_52,
       rd_hit_oh_0_51,
       rd_hit_oh_0_50,
       rd_hit_oh_0_49,
       rd_hit_oh_0_48,
       rd_hit_oh_0_47,
       rd_hit_oh_0_46,
       rd_hit_oh_0_45,
       rd_hit_oh_0_44,
       rd_hit_oh_0_43,
       rd_hit_oh_0_42,
       rd_hit_oh_0_41,
       rd_hit_oh_0_40,
       rd_hit_oh_0_39,
       rd_hit_oh_0_38,
       rd_hit_oh_0_37,
       rd_hit_oh_0_36,
       rd_hit_oh_0_35,
       rd_hit_oh_0_34,
       rd_hit_oh_0_33,
       crat_32_valid & crat_32_lr == io_rd_0},
     |(_io_pprd_0_T_1073[30:15]),
     |(_io_pprd_0_T_1075[14:7]),
     |(_io_pprd_0_T_1077[6:3]),
     |(_io_pprd_0_T_1079[2:1]),
     _io_pprd_0_T_1079[2] | _io_pprd_0_T_1079[0]};
  wire        rj_hit_oh_1_33 = crat_33_valid & crat_33_lr == io_rj_1;
  wire        rk_hit_oh_1_33 = crat_33_valid & crat_33_lr == io_rk_1;
  wire        rd_hit_oh_1_33 = crat_33_valid & crat_33_lr == io_rd_1;
  wire        rj_hit_oh_1_34 = crat_34_valid & crat_34_lr == io_rj_1;
  wire        rk_hit_oh_1_34 = crat_34_valid & crat_34_lr == io_rk_1;
  wire        rd_hit_oh_1_34 = crat_34_valid & crat_34_lr == io_rd_1;
  wire        rj_hit_oh_1_35 = crat_35_valid & crat_35_lr == io_rj_1;
  wire        rk_hit_oh_1_35 = crat_35_valid & crat_35_lr == io_rk_1;
  wire        rd_hit_oh_1_35 = crat_35_valid & crat_35_lr == io_rd_1;
  wire        rj_hit_oh_1_36 = crat_36_valid & crat_36_lr == io_rj_1;
  wire        rk_hit_oh_1_36 = crat_36_valid & crat_36_lr == io_rk_1;
  wire        rd_hit_oh_1_36 = crat_36_valid & crat_36_lr == io_rd_1;
  wire        rj_hit_oh_1_37 = crat_37_valid & crat_37_lr == io_rj_1;
  wire        rk_hit_oh_1_37 = crat_37_valid & crat_37_lr == io_rk_1;
  wire        rd_hit_oh_1_37 = crat_37_valid & crat_37_lr == io_rd_1;
  wire        rj_hit_oh_1_38 = crat_38_valid & crat_38_lr == io_rj_1;
  wire        rk_hit_oh_1_38 = crat_38_valid & crat_38_lr == io_rk_1;
  wire        rd_hit_oh_1_38 = crat_38_valid & crat_38_lr == io_rd_1;
  wire        rj_hit_oh_1_39 = crat_39_valid & crat_39_lr == io_rj_1;
  wire        rk_hit_oh_1_39 = crat_39_valid & crat_39_lr == io_rk_1;
  wire        rd_hit_oh_1_39 = crat_39_valid & crat_39_lr == io_rd_1;
  wire        rj_hit_oh_1_40 = crat_40_valid & crat_40_lr == io_rj_1;
  wire        rk_hit_oh_1_40 = crat_40_valid & crat_40_lr == io_rk_1;
  wire        rd_hit_oh_1_40 = crat_40_valid & crat_40_lr == io_rd_1;
  wire        rj_hit_oh_1_41 = crat_41_valid & crat_41_lr == io_rj_1;
  wire        rk_hit_oh_1_41 = crat_41_valid & crat_41_lr == io_rk_1;
  wire        rd_hit_oh_1_41 = crat_41_valid & crat_41_lr == io_rd_1;
  wire        rj_hit_oh_1_42 = crat_42_valid & crat_42_lr == io_rj_1;
  wire        rk_hit_oh_1_42 = crat_42_valid & crat_42_lr == io_rk_1;
  wire        rd_hit_oh_1_42 = crat_42_valid & crat_42_lr == io_rd_1;
  wire        rj_hit_oh_1_43 = crat_43_valid & crat_43_lr == io_rj_1;
  wire        rk_hit_oh_1_43 = crat_43_valid & crat_43_lr == io_rk_1;
  wire        rd_hit_oh_1_43 = crat_43_valid & crat_43_lr == io_rd_1;
  wire        rj_hit_oh_1_44 = crat_44_valid & crat_44_lr == io_rj_1;
  wire        rk_hit_oh_1_44 = crat_44_valid & crat_44_lr == io_rk_1;
  wire        rd_hit_oh_1_44 = crat_44_valid & crat_44_lr == io_rd_1;
  wire        rj_hit_oh_1_45 = crat_45_valid & crat_45_lr == io_rj_1;
  wire        rk_hit_oh_1_45 = crat_45_valid & crat_45_lr == io_rk_1;
  wire        rd_hit_oh_1_45 = crat_45_valid & crat_45_lr == io_rd_1;
  wire        rj_hit_oh_1_46 = crat_46_valid & crat_46_lr == io_rj_1;
  wire        rk_hit_oh_1_46 = crat_46_valid & crat_46_lr == io_rk_1;
  wire        rd_hit_oh_1_46 = crat_46_valid & crat_46_lr == io_rd_1;
  wire        rj_hit_oh_1_47 = crat_47_valid & crat_47_lr == io_rj_1;
  wire        rk_hit_oh_1_47 = crat_47_valid & crat_47_lr == io_rk_1;
  wire        rd_hit_oh_1_47 = crat_47_valid & crat_47_lr == io_rd_1;
  wire        rj_hit_oh_1_48 = crat_48_valid & crat_48_lr == io_rj_1;
  wire        rk_hit_oh_1_48 = crat_48_valid & crat_48_lr == io_rk_1;
  wire        rd_hit_oh_1_48 = crat_48_valid & crat_48_lr == io_rd_1;
  wire        rj_hit_oh_1_49 = crat_49_valid & crat_49_lr == io_rj_1;
  wire        rk_hit_oh_1_49 = crat_49_valid & crat_49_lr == io_rk_1;
  wire        rd_hit_oh_1_49 = crat_49_valid & crat_49_lr == io_rd_1;
  wire        rj_hit_oh_1_50 = crat_50_valid & crat_50_lr == io_rj_1;
  wire        rk_hit_oh_1_50 = crat_50_valid & crat_50_lr == io_rk_1;
  wire        rd_hit_oh_1_50 = crat_50_valid & crat_50_lr == io_rd_1;
  wire        rj_hit_oh_1_51 = crat_51_valid & crat_51_lr == io_rj_1;
  wire        rk_hit_oh_1_51 = crat_51_valid & crat_51_lr == io_rk_1;
  wire        rd_hit_oh_1_51 = crat_51_valid & crat_51_lr == io_rd_1;
  wire        rj_hit_oh_1_52 = crat_52_valid & crat_52_lr == io_rj_1;
  wire        rk_hit_oh_1_52 = crat_52_valid & crat_52_lr == io_rk_1;
  wire        rd_hit_oh_1_52 = crat_52_valid & crat_52_lr == io_rd_1;
  wire        rj_hit_oh_1_53 = crat_53_valid & crat_53_lr == io_rj_1;
  wire        rk_hit_oh_1_53 = crat_53_valid & crat_53_lr == io_rk_1;
  wire        rd_hit_oh_1_53 = crat_53_valid & crat_53_lr == io_rd_1;
  wire        rj_hit_oh_1_54 = crat_54_valid & crat_54_lr == io_rj_1;
  wire        rk_hit_oh_1_54 = crat_54_valid & crat_54_lr == io_rk_1;
  wire        rd_hit_oh_1_54 = crat_54_valid & crat_54_lr == io_rd_1;
  wire        rj_hit_oh_1_55 = crat_55_valid & crat_55_lr == io_rj_1;
  wire        rk_hit_oh_1_55 = crat_55_valid & crat_55_lr == io_rk_1;
  wire        rd_hit_oh_1_55 = crat_55_valid & crat_55_lr == io_rd_1;
  wire        rj_hit_oh_1_56 = crat_56_valid & crat_56_lr == io_rj_1;
  wire        rk_hit_oh_1_56 = crat_56_valid & crat_56_lr == io_rk_1;
  wire        rd_hit_oh_1_56 = crat_56_valid & crat_56_lr == io_rd_1;
  wire        rj_hit_oh_1_57 = crat_57_valid & crat_57_lr == io_rj_1;
  wire        rk_hit_oh_1_57 = crat_57_valid & crat_57_lr == io_rk_1;
  wire        rd_hit_oh_1_57 = crat_57_valid & crat_57_lr == io_rd_1;
  wire        rj_hit_oh_1_58 = crat_58_valid & crat_58_lr == io_rj_1;
  wire        rk_hit_oh_1_58 = crat_58_valid & crat_58_lr == io_rk_1;
  wire        rd_hit_oh_1_58 = crat_58_valid & crat_58_lr == io_rd_1;
  wire        rj_hit_oh_1_59 = crat_59_valid & crat_59_lr == io_rj_1;
  wire        rk_hit_oh_1_59 = crat_59_valid & crat_59_lr == io_rk_1;
  wire        rd_hit_oh_1_59 = crat_59_valid & crat_59_lr == io_rd_1;
  wire        rj_hit_oh_1_60 = crat_60_valid & crat_60_lr == io_rj_1;
  wire        rk_hit_oh_1_60 = crat_60_valid & crat_60_lr == io_rk_1;
  wire        rd_hit_oh_1_60 = crat_60_valid & crat_60_lr == io_rd_1;
  wire        rj_hit_oh_1_61 = crat_61_valid & crat_61_lr == io_rj_1;
  wire        rk_hit_oh_1_61 = crat_61_valid & crat_61_lr == io_rk_1;
  wire        rd_hit_oh_1_61 = crat_61_valid & crat_61_lr == io_rd_1;
  wire        rj_hit_oh_1_62 = crat_62_valid & crat_62_lr == io_rj_1;
  wire        rk_hit_oh_1_62 = crat_62_valid & crat_62_lr == io_rk_1;
  wire        rd_hit_oh_1_62 = crat_62_valid & crat_62_lr == io_rd_1;
  wire        rj_hit_oh_1_63 = crat_63_valid & crat_63_lr == io_rj_1;
  wire        rk_hit_oh_1_63 = crat_63_valid & crat_63_lr == io_rk_1;
  wire        rd_hit_oh_1_63 = crat_63_valid & crat_63_lr == io_rd_1;
  wire [30:0] _io_prj_1_T_1073 =
    {rj_hit_oh_1_63,
     rj_hit_oh_1_62,
     rj_hit_oh_1_61,
     rj_hit_oh_1_60,
     rj_hit_oh_1_59,
     rj_hit_oh_1_58,
     rj_hit_oh_1_57,
     rj_hit_oh_1_56,
     rj_hit_oh_1_55,
     rj_hit_oh_1_54,
     rj_hit_oh_1_53,
     rj_hit_oh_1_52,
     rj_hit_oh_1_51,
     rj_hit_oh_1_50,
     rj_hit_oh_1_49,
     rj_hit_oh_1_48,
     rj_hit_oh_1_47,
     rj_hit_oh_1_46,
     rj_hit_oh_1_45,
     rj_hit_oh_1_44,
     rj_hit_oh_1_43,
     rj_hit_oh_1_42,
     rj_hit_oh_1_41,
     rj_hit_oh_1_40,
     rj_hit_oh_1_39,
     rj_hit_oh_1_38,
     rj_hit_oh_1_37,
     rj_hit_oh_1_36,
     rj_hit_oh_1_35,
     rj_hit_oh_1_34,
     rj_hit_oh_1_33}
    | {crat_31_valid & crat_31_lr == io_rj_1,
       crat_30_valid & crat_30_lr == io_rj_1,
       crat_29_valid & crat_29_lr == io_rj_1,
       crat_28_valid & crat_28_lr == io_rj_1,
       crat_27_valid & crat_27_lr == io_rj_1,
       crat_26_valid & crat_26_lr == io_rj_1,
       crat_25_valid & crat_25_lr == io_rj_1,
       crat_24_valid & crat_24_lr == io_rj_1,
       crat_23_valid & crat_23_lr == io_rj_1,
       crat_22_valid & crat_22_lr == io_rj_1,
       crat_21_valid & crat_21_lr == io_rj_1,
       crat_20_valid & crat_20_lr == io_rj_1,
       crat_19_valid & crat_19_lr == io_rj_1,
       crat_18_valid & crat_18_lr == io_rj_1,
       crat_17_valid & crat_17_lr == io_rj_1,
       crat_16_valid & crat_16_lr == io_rj_1,
       crat_15_valid & crat_15_lr == io_rj_1,
       crat_14_valid & crat_14_lr == io_rj_1,
       crat_13_valid & crat_13_lr == io_rj_1,
       crat_12_valid & crat_12_lr == io_rj_1,
       crat_11_valid & crat_11_lr == io_rj_1,
       crat_10_valid & crat_10_lr == io_rj_1,
       crat_9_valid & crat_9_lr == io_rj_1,
       crat_8_valid & crat_8_lr == io_rj_1,
       crat_7_valid & crat_7_lr == io_rj_1,
       crat_6_valid & crat_6_lr == io_rj_1,
       crat_5_valid & crat_5_lr == io_rj_1,
       crat_4_valid & crat_4_lr == io_rj_1,
       crat_3_valid & crat_3_lr == io_rj_1,
       crat_2_valid & crat_2_lr == io_rj_1,
       crat_1_valid & crat_1_lr == io_rj_1};
  wire [14:0] _io_prj_1_T_1075 = _io_prj_1_T_1073[30:16] | _io_prj_1_T_1073[14:0];
  wire [6:0]  _io_prj_1_T_1077 = _io_prj_1_T_1075[14:8] | _io_prj_1_T_1075[6:0];
  wire [2:0]  _io_prj_1_T_1079 = _io_prj_1_T_1077[6:4] | _io_prj_1_T_1077[2:0];
  wire [30:0] _io_prk_1_T_1073 =
    {rk_hit_oh_1_63,
     rk_hit_oh_1_62,
     rk_hit_oh_1_61,
     rk_hit_oh_1_60,
     rk_hit_oh_1_59,
     rk_hit_oh_1_58,
     rk_hit_oh_1_57,
     rk_hit_oh_1_56,
     rk_hit_oh_1_55,
     rk_hit_oh_1_54,
     rk_hit_oh_1_53,
     rk_hit_oh_1_52,
     rk_hit_oh_1_51,
     rk_hit_oh_1_50,
     rk_hit_oh_1_49,
     rk_hit_oh_1_48,
     rk_hit_oh_1_47,
     rk_hit_oh_1_46,
     rk_hit_oh_1_45,
     rk_hit_oh_1_44,
     rk_hit_oh_1_43,
     rk_hit_oh_1_42,
     rk_hit_oh_1_41,
     rk_hit_oh_1_40,
     rk_hit_oh_1_39,
     rk_hit_oh_1_38,
     rk_hit_oh_1_37,
     rk_hit_oh_1_36,
     rk_hit_oh_1_35,
     rk_hit_oh_1_34,
     rk_hit_oh_1_33}
    | {crat_31_valid & crat_31_lr == io_rk_1,
       crat_30_valid & crat_30_lr == io_rk_1,
       crat_29_valid & crat_29_lr == io_rk_1,
       crat_28_valid & crat_28_lr == io_rk_1,
       crat_27_valid & crat_27_lr == io_rk_1,
       crat_26_valid & crat_26_lr == io_rk_1,
       crat_25_valid & crat_25_lr == io_rk_1,
       crat_24_valid & crat_24_lr == io_rk_1,
       crat_23_valid & crat_23_lr == io_rk_1,
       crat_22_valid & crat_22_lr == io_rk_1,
       crat_21_valid & crat_21_lr == io_rk_1,
       crat_20_valid & crat_20_lr == io_rk_1,
       crat_19_valid & crat_19_lr == io_rk_1,
       crat_18_valid & crat_18_lr == io_rk_1,
       crat_17_valid & crat_17_lr == io_rk_1,
       crat_16_valid & crat_16_lr == io_rk_1,
       crat_15_valid & crat_15_lr == io_rk_1,
       crat_14_valid & crat_14_lr == io_rk_1,
       crat_13_valid & crat_13_lr == io_rk_1,
       crat_12_valid & crat_12_lr == io_rk_1,
       crat_11_valid & crat_11_lr == io_rk_1,
       crat_10_valid & crat_10_lr == io_rk_1,
       crat_9_valid & crat_9_lr == io_rk_1,
       crat_8_valid & crat_8_lr == io_rk_1,
       crat_7_valid & crat_7_lr == io_rk_1,
       crat_6_valid & crat_6_lr == io_rk_1,
       crat_5_valid & crat_5_lr == io_rk_1,
       crat_4_valid & crat_4_lr == io_rk_1,
       crat_3_valid & crat_3_lr == io_rk_1,
       crat_2_valid & crat_2_lr == io_rk_1,
       crat_1_valid & crat_1_lr == io_rk_1};
  wire [14:0] _io_prk_1_T_1075 = _io_prk_1_T_1073[30:16] | _io_prk_1_T_1073[14:0];
  wire [6:0]  _io_prk_1_T_1077 = _io_prk_1_T_1075[14:8] | _io_prk_1_T_1075[6:0];
  wire [2:0]  _io_prk_1_T_1079 = _io_prk_1_T_1077[6:4] | _io_prk_1_T_1077[2:0];
  wire [30:0] _io_pprd_1_T_1073 =
    {rd_hit_oh_1_63,
     rd_hit_oh_1_62,
     rd_hit_oh_1_61,
     rd_hit_oh_1_60,
     rd_hit_oh_1_59,
     rd_hit_oh_1_58,
     rd_hit_oh_1_57,
     rd_hit_oh_1_56,
     rd_hit_oh_1_55,
     rd_hit_oh_1_54,
     rd_hit_oh_1_53,
     rd_hit_oh_1_52,
     rd_hit_oh_1_51,
     rd_hit_oh_1_50,
     rd_hit_oh_1_49,
     rd_hit_oh_1_48,
     rd_hit_oh_1_47,
     rd_hit_oh_1_46,
     rd_hit_oh_1_45,
     rd_hit_oh_1_44,
     rd_hit_oh_1_43,
     rd_hit_oh_1_42,
     rd_hit_oh_1_41,
     rd_hit_oh_1_40,
     rd_hit_oh_1_39,
     rd_hit_oh_1_38,
     rd_hit_oh_1_37,
     rd_hit_oh_1_36,
     rd_hit_oh_1_35,
     rd_hit_oh_1_34,
     rd_hit_oh_1_33}
    | {crat_31_valid & crat_31_lr == io_rd_1,
       crat_30_valid & crat_30_lr == io_rd_1,
       crat_29_valid & crat_29_lr == io_rd_1,
       crat_28_valid & crat_28_lr == io_rd_1,
       crat_27_valid & crat_27_lr == io_rd_1,
       crat_26_valid & crat_26_lr == io_rd_1,
       crat_25_valid & crat_25_lr == io_rd_1,
       crat_24_valid & crat_24_lr == io_rd_1,
       crat_23_valid & crat_23_lr == io_rd_1,
       crat_22_valid & crat_22_lr == io_rd_1,
       crat_21_valid & crat_21_lr == io_rd_1,
       crat_20_valid & crat_20_lr == io_rd_1,
       crat_19_valid & crat_19_lr == io_rd_1,
       crat_18_valid & crat_18_lr == io_rd_1,
       crat_17_valid & crat_17_lr == io_rd_1,
       crat_16_valid & crat_16_lr == io_rd_1,
       crat_15_valid & crat_15_lr == io_rd_1,
       crat_14_valid & crat_14_lr == io_rd_1,
       crat_13_valid & crat_13_lr == io_rd_1,
       crat_12_valid & crat_12_lr == io_rd_1,
       crat_11_valid & crat_11_lr == io_rd_1,
       crat_10_valid & crat_10_lr == io_rd_1,
       crat_9_valid & crat_9_lr == io_rd_1,
       crat_8_valid & crat_8_lr == io_rd_1,
       crat_7_valid & crat_7_lr == io_rd_1,
       crat_6_valid & crat_6_lr == io_rd_1,
       crat_5_valid & crat_5_lr == io_rd_1,
       crat_4_valid & crat_4_lr == io_rd_1,
       crat_3_valid & crat_3_lr == io_rd_1,
       crat_2_valid & crat_2_lr == io_rd_1,
       crat_1_valid & crat_1_lr == io_rd_1};
  wire [14:0] _io_pprd_1_T_1075 = _io_pprd_1_T_1073[30:16] | _io_pprd_1_T_1073[14:0];
  wire [6:0]  _io_pprd_1_T_1077 = _io_pprd_1_T_1075[14:8] | _io_pprd_1_T_1075[6:0];
  wire [2:0]  _io_pprd_1_T_1079 = _io_pprd_1_T_1077[6:4] | _io_pprd_1_T_1077[2:0];
  wire [5:0]  _io_pprd_1_output =
    {|{rd_hit_oh_1_63,
       rd_hit_oh_1_62,
       rd_hit_oh_1_61,
       rd_hit_oh_1_60,
       rd_hit_oh_1_59,
       rd_hit_oh_1_58,
       rd_hit_oh_1_57,
       rd_hit_oh_1_56,
       rd_hit_oh_1_55,
       rd_hit_oh_1_54,
       rd_hit_oh_1_53,
       rd_hit_oh_1_52,
       rd_hit_oh_1_51,
       rd_hit_oh_1_50,
       rd_hit_oh_1_49,
       rd_hit_oh_1_48,
       rd_hit_oh_1_47,
       rd_hit_oh_1_46,
       rd_hit_oh_1_45,
       rd_hit_oh_1_44,
       rd_hit_oh_1_43,
       rd_hit_oh_1_42,
       rd_hit_oh_1_41,
       rd_hit_oh_1_40,
       rd_hit_oh_1_39,
       rd_hit_oh_1_38,
       rd_hit_oh_1_37,
       rd_hit_oh_1_36,
       rd_hit_oh_1_35,
       rd_hit_oh_1_34,
       rd_hit_oh_1_33,
       crat_32_valid & crat_32_lr == io_rd_1},
     |(_io_pprd_1_T_1073[30:15]),
     |(_io_pprd_1_T_1075[14:7]),
     |(_io_pprd_1_T_1077[6:3]),
     |(_io_pprd_1_T_1079[2:1]),
     _io_pprd_1_T_1079[2] | _io_pprd_1_T_1079[0]};
  wire        rj_hit_oh_2_33 = crat_33_valid & crat_33_lr == io_rj_2;
  wire        rk_hit_oh_2_33 = crat_33_valid & crat_33_lr == io_rk_2;
  wire        rd_hit_oh_2_33 = crat_33_valid & crat_33_lr == io_rd_2;
  wire        rj_hit_oh_2_34 = crat_34_valid & crat_34_lr == io_rj_2;
  wire        rk_hit_oh_2_34 = crat_34_valid & crat_34_lr == io_rk_2;
  wire        rd_hit_oh_2_34 = crat_34_valid & crat_34_lr == io_rd_2;
  wire        rj_hit_oh_2_35 = crat_35_valid & crat_35_lr == io_rj_2;
  wire        rk_hit_oh_2_35 = crat_35_valid & crat_35_lr == io_rk_2;
  wire        rd_hit_oh_2_35 = crat_35_valid & crat_35_lr == io_rd_2;
  wire        rj_hit_oh_2_36 = crat_36_valid & crat_36_lr == io_rj_2;
  wire        rk_hit_oh_2_36 = crat_36_valid & crat_36_lr == io_rk_2;
  wire        rd_hit_oh_2_36 = crat_36_valid & crat_36_lr == io_rd_2;
  wire        rj_hit_oh_2_37 = crat_37_valid & crat_37_lr == io_rj_2;
  wire        rk_hit_oh_2_37 = crat_37_valid & crat_37_lr == io_rk_2;
  wire        rd_hit_oh_2_37 = crat_37_valid & crat_37_lr == io_rd_2;
  wire        rj_hit_oh_2_38 = crat_38_valid & crat_38_lr == io_rj_2;
  wire        rk_hit_oh_2_38 = crat_38_valid & crat_38_lr == io_rk_2;
  wire        rd_hit_oh_2_38 = crat_38_valid & crat_38_lr == io_rd_2;
  wire        rj_hit_oh_2_39 = crat_39_valid & crat_39_lr == io_rj_2;
  wire        rk_hit_oh_2_39 = crat_39_valid & crat_39_lr == io_rk_2;
  wire        rd_hit_oh_2_39 = crat_39_valid & crat_39_lr == io_rd_2;
  wire        rj_hit_oh_2_40 = crat_40_valid & crat_40_lr == io_rj_2;
  wire        rk_hit_oh_2_40 = crat_40_valid & crat_40_lr == io_rk_2;
  wire        rd_hit_oh_2_40 = crat_40_valid & crat_40_lr == io_rd_2;
  wire        rj_hit_oh_2_41 = crat_41_valid & crat_41_lr == io_rj_2;
  wire        rk_hit_oh_2_41 = crat_41_valid & crat_41_lr == io_rk_2;
  wire        rd_hit_oh_2_41 = crat_41_valid & crat_41_lr == io_rd_2;
  wire        rj_hit_oh_2_42 = crat_42_valid & crat_42_lr == io_rj_2;
  wire        rk_hit_oh_2_42 = crat_42_valid & crat_42_lr == io_rk_2;
  wire        rd_hit_oh_2_42 = crat_42_valid & crat_42_lr == io_rd_2;
  wire        rj_hit_oh_2_43 = crat_43_valid & crat_43_lr == io_rj_2;
  wire        rk_hit_oh_2_43 = crat_43_valid & crat_43_lr == io_rk_2;
  wire        rd_hit_oh_2_43 = crat_43_valid & crat_43_lr == io_rd_2;
  wire        rj_hit_oh_2_44 = crat_44_valid & crat_44_lr == io_rj_2;
  wire        rk_hit_oh_2_44 = crat_44_valid & crat_44_lr == io_rk_2;
  wire        rd_hit_oh_2_44 = crat_44_valid & crat_44_lr == io_rd_2;
  wire        rj_hit_oh_2_45 = crat_45_valid & crat_45_lr == io_rj_2;
  wire        rk_hit_oh_2_45 = crat_45_valid & crat_45_lr == io_rk_2;
  wire        rd_hit_oh_2_45 = crat_45_valid & crat_45_lr == io_rd_2;
  wire        rj_hit_oh_2_46 = crat_46_valid & crat_46_lr == io_rj_2;
  wire        rk_hit_oh_2_46 = crat_46_valid & crat_46_lr == io_rk_2;
  wire        rd_hit_oh_2_46 = crat_46_valid & crat_46_lr == io_rd_2;
  wire        rj_hit_oh_2_47 = crat_47_valid & crat_47_lr == io_rj_2;
  wire        rk_hit_oh_2_47 = crat_47_valid & crat_47_lr == io_rk_2;
  wire        rd_hit_oh_2_47 = crat_47_valid & crat_47_lr == io_rd_2;
  wire        rj_hit_oh_2_48 = crat_48_valid & crat_48_lr == io_rj_2;
  wire        rk_hit_oh_2_48 = crat_48_valid & crat_48_lr == io_rk_2;
  wire        rd_hit_oh_2_48 = crat_48_valid & crat_48_lr == io_rd_2;
  wire        rj_hit_oh_2_49 = crat_49_valid & crat_49_lr == io_rj_2;
  wire        rk_hit_oh_2_49 = crat_49_valid & crat_49_lr == io_rk_2;
  wire        rd_hit_oh_2_49 = crat_49_valid & crat_49_lr == io_rd_2;
  wire        rj_hit_oh_2_50 = crat_50_valid & crat_50_lr == io_rj_2;
  wire        rk_hit_oh_2_50 = crat_50_valid & crat_50_lr == io_rk_2;
  wire        rd_hit_oh_2_50 = crat_50_valid & crat_50_lr == io_rd_2;
  wire        rj_hit_oh_2_51 = crat_51_valid & crat_51_lr == io_rj_2;
  wire        rk_hit_oh_2_51 = crat_51_valid & crat_51_lr == io_rk_2;
  wire        rd_hit_oh_2_51 = crat_51_valid & crat_51_lr == io_rd_2;
  wire        rj_hit_oh_2_52 = crat_52_valid & crat_52_lr == io_rj_2;
  wire        rk_hit_oh_2_52 = crat_52_valid & crat_52_lr == io_rk_2;
  wire        rd_hit_oh_2_52 = crat_52_valid & crat_52_lr == io_rd_2;
  wire        rj_hit_oh_2_53 = crat_53_valid & crat_53_lr == io_rj_2;
  wire        rk_hit_oh_2_53 = crat_53_valid & crat_53_lr == io_rk_2;
  wire        rd_hit_oh_2_53 = crat_53_valid & crat_53_lr == io_rd_2;
  wire        rj_hit_oh_2_54 = crat_54_valid & crat_54_lr == io_rj_2;
  wire        rk_hit_oh_2_54 = crat_54_valid & crat_54_lr == io_rk_2;
  wire        rd_hit_oh_2_54 = crat_54_valid & crat_54_lr == io_rd_2;
  wire        rj_hit_oh_2_55 = crat_55_valid & crat_55_lr == io_rj_2;
  wire        rk_hit_oh_2_55 = crat_55_valid & crat_55_lr == io_rk_2;
  wire        rd_hit_oh_2_55 = crat_55_valid & crat_55_lr == io_rd_2;
  wire        rj_hit_oh_2_56 = crat_56_valid & crat_56_lr == io_rj_2;
  wire        rk_hit_oh_2_56 = crat_56_valid & crat_56_lr == io_rk_2;
  wire        rd_hit_oh_2_56 = crat_56_valid & crat_56_lr == io_rd_2;
  wire        rj_hit_oh_2_57 = crat_57_valid & crat_57_lr == io_rj_2;
  wire        rk_hit_oh_2_57 = crat_57_valid & crat_57_lr == io_rk_2;
  wire        rd_hit_oh_2_57 = crat_57_valid & crat_57_lr == io_rd_2;
  wire        rj_hit_oh_2_58 = crat_58_valid & crat_58_lr == io_rj_2;
  wire        rk_hit_oh_2_58 = crat_58_valid & crat_58_lr == io_rk_2;
  wire        rd_hit_oh_2_58 = crat_58_valid & crat_58_lr == io_rd_2;
  wire        rj_hit_oh_2_59 = crat_59_valid & crat_59_lr == io_rj_2;
  wire        rk_hit_oh_2_59 = crat_59_valid & crat_59_lr == io_rk_2;
  wire        rd_hit_oh_2_59 = crat_59_valid & crat_59_lr == io_rd_2;
  wire        rj_hit_oh_2_60 = crat_60_valid & crat_60_lr == io_rj_2;
  wire        rk_hit_oh_2_60 = crat_60_valid & crat_60_lr == io_rk_2;
  wire        rd_hit_oh_2_60 = crat_60_valid & crat_60_lr == io_rd_2;
  wire        rj_hit_oh_2_61 = crat_61_valid & crat_61_lr == io_rj_2;
  wire        rk_hit_oh_2_61 = crat_61_valid & crat_61_lr == io_rk_2;
  wire        rd_hit_oh_2_61 = crat_61_valid & crat_61_lr == io_rd_2;
  wire        rj_hit_oh_2_62 = crat_62_valid & crat_62_lr == io_rj_2;
  wire        rk_hit_oh_2_62 = crat_62_valid & crat_62_lr == io_rk_2;
  wire        rd_hit_oh_2_62 = crat_62_valid & crat_62_lr == io_rd_2;
  wire        rj_hit_oh_2_63 = crat_63_valid & crat_63_lr == io_rj_2;
  wire        rk_hit_oh_2_63 = crat_63_valid & crat_63_lr == io_rk_2;
  wire        rd_hit_oh_2_63 = crat_63_valid & crat_63_lr == io_rd_2;
  wire [30:0] _io_prj_2_T_1073 =
    {rj_hit_oh_2_63,
     rj_hit_oh_2_62,
     rj_hit_oh_2_61,
     rj_hit_oh_2_60,
     rj_hit_oh_2_59,
     rj_hit_oh_2_58,
     rj_hit_oh_2_57,
     rj_hit_oh_2_56,
     rj_hit_oh_2_55,
     rj_hit_oh_2_54,
     rj_hit_oh_2_53,
     rj_hit_oh_2_52,
     rj_hit_oh_2_51,
     rj_hit_oh_2_50,
     rj_hit_oh_2_49,
     rj_hit_oh_2_48,
     rj_hit_oh_2_47,
     rj_hit_oh_2_46,
     rj_hit_oh_2_45,
     rj_hit_oh_2_44,
     rj_hit_oh_2_43,
     rj_hit_oh_2_42,
     rj_hit_oh_2_41,
     rj_hit_oh_2_40,
     rj_hit_oh_2_39,
     rj_hit_oh_2_38,
     rj_hit_oh_2_37,
     rj_hit_oh_2_36,
     rj_hit_oh_2_35,
     rj_hit_oh_2_34,
     rj_hit_oh_2_33}
    | {crat_31_valid & crat_31_lr == io_rj_2,
       crat_30_valid & crat_30_lr == io_rj_2,
       crat_29_valid & crat_29_lr == io_rj_2,
       crat_28_valid & crat_28_lr == io_rj_2,
       crat_27_valid & crat_27_lr == io_rj_2,
       crat_26_valid & crat_26_lr == io_rj_2,
       crat_25_valid & crat_25_lr == io_rj_2,
       crat_24_valid & crat_24_lr == io_rj_2,
       crat_23_valid & crat_23_lr == io_rj_2,
       crat_22_valid & crat_22_lr == io_rj_2,
       crat_21_valid & crat_21_lr == io_rj_2,
       crat_20_valid & crat_20_lr == io_rj_2,
       crat_19_valid & crat_19_lr == io_rj_2,
       crat_18_valid & crat_18_lr == io_rj_2,
       crat_17_valid & crat_17_lr == io_rj_2,
       crat_16_valid & crat_16_lr == io_rj_2,
       crat_15_valid & crat_15_lr == io_rj_2,
       crat_14_valid & crat_14_lr == io_rj_2,
       crat_13_valid & crat_13_lr == io_rj_2,
       crat_12_valid & crat_12_lr == io_rj_2,
       crat_11_valid & crat_11_lr == io_rj_2,
       crat_10_valid & crat_10_lr == io_rj_2,
       crat_9_valid & crat_9_lr == io_rj_2,
       crat_8_valid & crat_8_lr == io_rj_2,
       crat_7_valid & crat_7_lr == io_rj_2,
       crat_6_valid & crat_6_lr == io_rj_2,
       crat_5_valid & crat_5_lr == io_rj_2,
       crat_4_valid & crat_4_lr == io_rj_2,
       crat_3_valid & crat_3_lr == io_rj_2,
       crat_2_valid & crat_2_lr == io_rj_2,
       crat_1_valid & crat_1_lr == io_rj_2};
  wire [14:0] _io_prj_2_T_1075 = _io_prj_2_T_1073[30:16] | _io_prj_2_T_1073[14:0];
  wire [6:0]  _io_prj_2_T_1077 = _io_prj_2_T_1075[14:8] | _io_prj_2_T_1075[6:0];
  wire [2:0]  _io_prj_2_T_1079 = _io_prj_2_T_1077[6:4] | _io_prj_2_T_1077[2:0];
  wire [30:0] _io_prk_2_T_1073 =
    {rk_hit_oh_2_63,
     rk_hit_oh_2_62,
     rk_hit_oh_2_61,
     rk_hit_oh_2_60,
     rk_hit_oh_2_59,
     rk_hit_oh_2_58,
     rk_hit_oh_2_57,
     rk_hit_oh_2_56,
     rk_hit_oh_2_55,
     rk_hit_oh_2_54,
     rk_hit_oh_2_53,
     rk_hit_oh_2_52,
     rk_hit_oh_2_51,
     rk_hit_oh_2_50,
     rk_hit_oh_2_49,
     rk_hit_oh_2_48,
     rk_hit_oh_2_47,
     rk_hit_oh_2_46,
     rk_hit_oh_2_45,
     rk_hit_oh_2_44,
     rk_hit_oh_2_43,
     rk_hit_oh_2_42,
     rk_hit_oh_2_41,
     rk_hit_oh_2_40,
     rk_hit_oh_2_39,
     rk_hit_oh_2_38,
     rk_hit_oh_2_37,
     rk_hit_oh_2_36,
     rk_hit_oh_2_35,
     rk_hit_oh_2_34,
     rk_hit_oh_2_33}
    | {crat_31_valid & crat_31_lr == io_rk_2,
       crat_30_valid & crat_30_lr == io_rk_2,
       crat_29_valid & crat_29_lr == io_rk_2,
       crat_28_valid & crat_28_lr == io_rk_2,
       crat_27_valid & crat_27_lr == io_rk_2,
       crat_26_valid & crat_26_lr == io_rk_2,
       crat_25_valid & crat_25_lr == io_rk_2,
       crat_24_valid & crat_24_lr == io_rk_2,
       crat_23_valid & crat_23_lr == io_rk_2,
       crat_22_valid & crat_22_lr == io_rk_2,
       crat_21_valid & crat_21_lr == io_rk_2,
       crat_20_valid & crat_20_lr == io_rk_2,
       crat_19_valid & crat_19_lr == io_rk_2,
       crat_18_valid & crat_18_lr == io_rk_2,
       crat_17_valid & crat_17_lr == io_rk_2,
       crat_16_valid & crat_16_lr == io_rk_2,
       crat_15_valid & crat_15_lr == io_rk_2,
       crat_14_valid & crat_14_lr == io_rk_2,
       crat_13_valid & crat_13_lr == io_rk_2,
       crat_12_valid & crat_12_lr == io_rk_2,
       crat_11_valid & crat_11_lr == io_rk_2,
       crat_10_valid & crat_10_lr == io_rk_2,
       crat_9_valid & crat_9_lr == io_rk_2,
       crat_8_valid & crat_8_lr == io_rk_2,
       crat_7_valid & crat_7_lr == io_rk_2,
       crat_6_valid & crat_6_lr == io_rk_2,
       crat_5_valid & crat_5_lr == io_rk_2,
       crat_4_valid & crat_4_lr == io_rk_2,
       crat_3_valid & crat_3_lr == io_rk_2,
       crat_2_valid & crat_2_lr == io_rk_2,
       crat_1_valid & crat_1_lr == io_rk_2};
  wire [14:0] _io_prk_2_T_1075 = _io_prk_2_T_1073[30:16] | _io_prk_2_T_1073[14:0];
  wire [6:0]  _io_prk_2_T_1077 = _io_prk_2_T_1075[14:8] | _io_prk_2_T_1075[6:0];
  wire [2:0]  _io_prk_2_T_1079 = _io_prk_2_T_1077[6:4] | _io_prk_2_T_1077[2:0];
  wire [30:0] _io_pprd_2_T_1073 =
    {rd_hit_oh_2_63,
     rd_hit_oh_2_62,
     rd_hit_oh_2_61,
     rd_hit_oh_2_60,
     rd_hit_oh_2_59,
     rd_hit_oh_2_58,
     rd_hit_oh_2_57,
     rd_hit_oh_2_56,
     rd_hit_oh_2_55,
     rd_hit_oh_2_54,
     rd_hit_oh_2_53,
     rd_hit_oh_2_52,
     rd_hit_oh_2_51,
     rd_hit_oh_2_50,
     rd_hit_oh_2_49,
     rd_hit_oh_2_48,
     rd_hit_oh_2_47,
     rd_hit_oh_2_46,
     rd_hit_oh_2_45,
     rd_hit_oh_2_44,
     rd_hit_oh_2_43,
     rd_hit_oh_2_42,
     rd_hit_oh_2_41,
     rd_hit_oh_2_40,
     rd_hit_oh_2_39,
     rd_hit_oh_2_38,
     rd_hit_oh_2_37,
     rd_hit_oh_2_36,
     rd_hit_oh_2_35,
     rd_hit_oh_2_34,
     rd_hit_oh_2_33}
    | {crat_31_valid & crat_31_lr == io_rd_2,
       crat_30_valid & crat_30_lr == io_rd_2,
       crat_29_valid & crat_29_lr == io_rd_2,
       crat_28_valid & crat_28_lr == io_rd_2,
       crat_27_valid & crat_27_lr == io_rd_2,
       crat_26_valid & crat_26_lr == io_rd_2,
       crat_25_valid & crat_25_lr == io_rd_2,
       crat_24_valid & crat_24_lr == io_rd_2,
       crat_23_valid & crat_23_lr == io_rd_2,
       crat_22_valid & crat_22_lr == io_rd_2,
       crat_21_valid & crat_21_lr == io_rd_2,
       crat_20_valid & crat_20_lr == io_rd_2,
       crat_19_valid & crat_19_lr == io_rd_2,
       crat_18_valid & crat_18_lr == io_rd_2,
       crat_17_valid & crat_17_lr == io_rd_2,
       crat_16_valid & crat_16_lr == io_rd_2,
       crat_15_valid & crat_15_lr == io_rd_2,
       crat_14_valid & crat_14_lr == io_rd_2,
       crat_13_valid & crat_13_lr == io_rd_2,
       crat_12_valid & crat_12_lr == io_rd_2,
       crat_11_valid & crat_11_lr == io_rd_2,
       crat_10_valid & crat_10_lr == io_rd_2,
       crat_9_valid & crat_9_lr == io_rd_2,
       crat_8_valid & crat_8_lr == io_rd_2,
       crat_7_valid & crat_7_lr == io_rd_2,
       crat_6_valid & crat_6_lr == io_rd_2,
       crat_5_valid & crat_5_lr == io_rd_2,
       crat_4_valid & crat_4_lr == io_rd_2,
       crat_3_valid & crat_3_lr == io_rd_2,
       crat_2_valid & crat_2_lr == io_rd_2,
       crat_1_valid & crat_1_lr == io_rd_2};
  wire [14:0] _io_pprd_2_T_1075 = _io_pprd_2_T_1073[30:16] | _io_pprd_2_T_1073[14:0];
  wire [6:0]  _io_pprd_2_T_1077 = _io_pprd_2_T_1075[14:8] | _io_pprd_2_T_1075[6:0];
  wire [2:0]  _io_pprd_2_T_1079 = _io_pprd_2_T_1077[6:4] | _io_pprd_2_T_1077[2:0];
  wire [5:0]  _io_pprd_2_output =
    {|{rd_hit_oh_2_63,
       rd_hit_oh_2_62,
       rd_hit_oh_2_61,
       rd_hit_oh_2_60,
       rd_hit_oh_2_59,
       rd_hit_oh_2_58,
       rd_hit_oh_2_57,
       rd_hit_oh_2_56,
       rd_hit_oh_2_55,
       rd_hit_oh_2_54,
       rd_hit_oh_2_53,
       rd_hit_oh_2_52,
       rd_hit_oh_2_51,
       rd_hit_oh_2_50,
       rd_hit_oh_2_49,
       rd_hit_oh_2_48,
       rd_hit_oh_2_47,
       rd_hit_oh_2_46,
       rd_hit_oh_2_45,
       rd_hit_oh_2_44,
       rd_hit_oh_2_43,
       rd_hit_oh_2_42,
       rd_hit_oh_2_41,
       rd_hit_oh_2_40,
       rd_hit_oh_2_39,
       rd_hit_oh_2_38,
       rd_hit_oh_2_37,
       rd_hit_oh_2_36,
       rd_hit_oh_2_35,
       rd_hit_oh_2_34,
       rd_hit_oh_2_33,
       crat_32_valid & crat_32_lr == io_rd_2},
     |(_io_pprd_2_T_1073[30:15]),
     |(_io_pprd_2_T_1075[14:7]),
     |(_io_pprd_2_T_1077[6:3]),
     |(_io_pprd_2_T_1079[2:1]),
     _io_pprd_2_T_1079[2] | _io_pprd_2_T_1079[0]};
  wire        rj_hit_oh_3_33 = crat_33_valid & crat_33_lr == io_rj_3;
  wire        rk_hit_oh_3_33 = crat_33_valid & crat_33_lr == io_rk_3;
  wire        rd_hit_oh_3_33 = crat_33_valid & crat_33_lr == io_rd_3;
  wire        rj_hit_oh_3_34 = crat_34_valid & crat_34_lr == io_rj_3;
  wire        rk_hit_oh_3_34 = crat_34_valid & crat_34_lr == io_rk_3;
  wire        rd_hit_oh_3_34 = crat_34_valid & crat_34_lr == io_rd_3;
  wire        rj_hit_oh_3_35 = crat_35_valid & crat_35_lr == io_rj_3;
  wire        rk_hit_oh_3_35 = crat_35_valid & crat_35_lr == io_rk_3;
  wire        rd_hit_oh_3_35 = crat_35_valid & crat_35_lr == io_rd_3;
  wire        rj_hit_oh_3_36 = crat_36_valid & crat_36_lr == io_rj_3;
  wire        rk_hit_oh_3_36 = crat_36_valid & crat_36_lr == io_rk_3;
  wire        rd_hit_oh_3_36 = crat_36_valid & crat_36_lr == io_rd_3;
  wire        rj_hit_oh_3_37 = crat_37_valid & crat_37_lr == io_rj_3;
  wire        rk_hit_oh_3_37 = crat_37_valid & crat_37_lr == io_rk_3;
  wire        rd_hit_oh_3_37 = crat_37_valid & crat_37_lr == io_rd_3;
  wire        rj_hit_oh_3_38 = crat_38_valid & crat_38_lr == io_rj_3;
  wire        rk_hit_oh_3_38 = crat_38_valid & crat_38_lr == io_rk_3;
  wire        rd_hit_oh_3_38 = crat_38_valid & crat_38_lr == io_rd_3;
  wire        rj_hit_oh_3_39 = crat_39_valid & crat_39_lr == io_rj_3;
  wire        rk_hit_oh_3_39 = crat_39_valid & crat_39_lr == io_rk_3;
  wire        rd_hit_oh_3_39 = crat_39_valid & crat_39_lr == io_rd_3;
  wire        rj_hit_oh_3_40 = crat_40_valid & crat_40_lr == io_rj_3;
  wire        rk_hit_oh_3_40 = crat_40_valid & crat_40_lr == io_rk_3;
  wire        rd_hit_oh_3_40 = crat_40_valid & crat_40_lr == io_rd_3;
  wire        rj_hit_oh_3_41 = crat_41_valid & crat_41_lr == io_rj_3;
  wire        rk_hit_oh_3_41 = crat_41_valid & crat_41_lr == io_rk_3;
  wire        rd_hit_oh_3_41 = crat_41_valid & crat_41_lr == io_rd_3;
  wire        rj_hit_oh_3_42 = crat_42_valid & crat_42_lr == io_rj_3;
  wire        rk_hit_oh_3_42 = crat_42_valid & crat_42_lr == io_rk_3;
  wire        rd_hit_oh_3_42 = crat_42_valid & crat_42_lr == io_rd_3;
  wire        rj_hit_oh_3_43 = crat_43_valid & crat_43_lr == io_rj_3;
  wire        rk_hit_oh_3_43 = crat_43_valid & crat_43_lr == io_rk_3;
  wire        rd_hit_oh_3_43 = crat_43_valid & crat_43_lr == io_rd_3;
  wire        rj_hit_oh_3_44 = crat_44_valid & crat_44_lr == io_rj_3;
  wire        rk_hit_oh_3_44 = crat_44_valid & crat_44_lr == io_rk_3;
  wire        rd_hit_oh_3_44 = crat_44_valid & crat_44_lr == io_rd_3;
  wire        rj_hit_oh_3_45 = crat_45_valid & crat_45_lr == io_rj_3;
  wire        rk_hit_oh_3_45 = crat_45_valid & crat_45_lr == io_rk_3;
  wire        rd_hit_oh_3_45 = crat_45_valid & crat_45_lr == io_rd_3;
  wire        rj_hit_oh_3_46 = crat_46_valid & crat_46_lr == io_rj_3;
  wire        rk_hit_oh_3_46 = crat_46_valid & crat_46_lr == io_rk_3;
  wire        rd_hit_oh_3_46 = crat_46_valid & crat_46_lr == io_rd_3;
  wire        rj_hit_oh_3_47 = crat_47_valid & crat_47_lr == io_rj_3;
  wire        rk_hit_oh_3_47 = crat_47_valid & crat_47_lr == io_rk_3;
  wire        rd_hit_oh_3_47 = crat_47_valid & crat_47_lr == io_rd_3;
  wire        rj_hit_oh_3_48 = crat_48_valid & crat_48_lr == io_rj_3;
  wire        rk_hit_oh_3_48 = crat_48_valid & crat_48_lr == io_rk_3;
  wire        rd_hit_oh_3_48 = crat_48_valid & crat_48_lr == io_rd_3;
  wire        rj_hit_oh_3_49 = crat_49_valid & crat_49_lr == io_rj_3;
  wire        rk_hit_oh_3_49 = crat_49_valid & crat_49_lr == io_rk_3;
  wire        rd_hit_oh_3_49 = crat_49_valid & crat_49_lr == io_rd_3;
  wire        rj_hit_oh_3_50 = crat_50_valid & crat_50_lr == io_rj_3;
  wire        rk_hit_oh_3_50 = crat_50_valid & crat_50_lr == io_rk_3;
  wire        rd_hit_oh_3_50 = crat_50_valid & crat_50_lr == io_rd_3;
  wire        rj_hit_oh_3_51 = crat_51_valid & crat_51_lr == io_rj_3;
  wire        rk_hit_oh_3_51 = crat_51_valid & crat_51_lr == io_rk_3;
  wire        rd_hit_oh_3_51 = crat_51_valid & crat_51_lr == io_rd_3;
  wire        rj_hit_oh_3_52 = crat_52_valid & crat_52_lr == io_rj_3;
  wire        rk_hit_oh_3_52 = crat_52_valid & crat_52_lr == io_rk_3;
  wire        rd_hit_oh_3_52 = crat_52_valid & crat_52_lr == io_rd_3;
  wire        rj_hit_oh_3_53 = crat_53_valid & crat_53_lr == io_rj_3;
  wire        rk_hit_oh_3_53 = crat_53_valid & crat_53_lr == io_rk_3;
  wire        rd_hit_oh_3_53 = crat_53_valid & crat_53_lr == io_rd_3;
  wire        rj_hit_oh_3_54 = crat_54_valid & crat_54_lr == io_rj_3;
  wire        rk_hit_oh_3_54 = crat_54_valid & crat_54_lr == io_rk_3;
  wire        rd_hit_oh_3_54 = crat_54_valid & crat_54_lr == io_rd_3;
  wire        rj_hit_oh_3_55 = crat_55_valid & crat_55_lr == io_rj_3;
  wire        rk_hit_oh_3_55 = crat_55_valid & crat_55_lr == io_rk_3;
  wire        rd_hit_oh_3_55 = crat_55_valid & crat_55_lr == io_rd_3;
  wire        rj_hit_oh_3_56 = crat_56_valid & crat_56_lr == io_rj_3;
  wire        rk_hit_oh_3_56 = crat_56_valid & crat_56_lr == io_rk_3;
  wire        rd_hit_oh_3_56 = crat_56_valid & crat_56_lr == io_rd_3;
  wire        rj_hit_oh_3_57 = crat_57_valid & crat_57_lr == io_rj_3;
  wire        rk_hit_oh_3_57 = crat_57_valid & crat_57_lr == io_rk_3;
  wire        rd_hit_oh_3_57 = crat_57_valid & crat_57_lr == io_rd_3;
  wire        rj_hit_oh_3_58 = crat_58_valid & crat_58_lr == io_rj_3;
  wire        rk_hit_oh_3_58 = crat_58_valid & crat_58_lr == io_rk_3;
  wire        rd_hit_oh_3_58 = crat_58_valid & crat_58_lr == io_rd_3;
  wire        rj_hit_oh_3_59 = crat_59_valid & crat_59_lr == io_rj_3;
  wire        rk_hit_oh_3_59 = crat_59_valid & crat_59_lr == io_rk_3;
  wire        rd_hit_oh_3_59 = crat_59_valid & crat_59_lr == io_rd_3;
  wire        rj_hit_oh_3_60 = crat_60_valid & crat_60_lr == io_rj_3;
  wire        rk_hit_oh_3_60 = crat_60_valid & crat_60_lr == io_rk_3;
  wire        rd_hit_oh_3_60 = crat_60_valid & crat_60_lr == io_rd_3;
  wire        rj_hit_oh_3_61 = crat_61_valid & crat_61_lr == io_rj_3;
  wire        rk_hit_oh_3_61 = crat_61_valid & crat_61_lr == io_rk_3;
  wire        rd_hit_oh_3_61 = crat_61_valid & crat_61_lr == io_rd_3;
  wire        rj_hit_oh_3_62 = crat_62_valid & crat_62_lr == io_rj_3;
  wire        rk_hit_oh_3_62 = crat_62_valid & crat_62_lr == io_rk_3;
  wire        rd_hit_oh_3_62 = crat_62_valid & crat_62_lr == io_rd_3;
  wire        rj_hit_oh_3_63 = crat_63_valid & crat_63_lr == io_rj_3;
  wire        rk_hit_oh_3_63 = crat_63_valid & crat_63_lr == io_rk_3;
  wire        rd_hit_oh_3_63 = crat_63_valid & crat_63_lr == io_rd_3;
  wire [30:0] _io_prj_3_T_1073 =
    {rj_hit_oh_3_63,
     rj_hit_oh_3_62,
     rj_hit_oh_3_61,
     rj_hit_oh_3_60,
     rj_hit_oh_3_59,
     rj_hit_oh_3_58,
     rj_hit_oh_3_57,
     rj_hit_oh_3_56,
     rj_hit_oh_3_55,
     rj_hit_oh_3_54,
     rj_hit_oh_3_53,
     rj_hit_oh_3_52,
     rj_hit_oh_3_51,
     rj_hit_oh_3_50,
     rj_hit_oh_3_49,
     rj_hit_oh_3_48,
     rj_hit_oh_3_47,
     rj_hit_oh_3_46,
     rj_hit_oh_3_45,
     rj_hit_oh_3_44,
     rj_hit_oh_3_43,
     rj_hit_oh_3_42,
     rj_hit_oh_3_41,
     rj_hit_oh_3_40,
     rj_hit_oh_3_39,
     rj_hit_oh_3_38,
     rj_hit_oh_3_37,
     rj_hit_oh_3_36,
     rj_hit_oh_3_35,
     rj_hit_oh_3_34,
     rj_hit_oh_3_33}
    | {crat_31_valid & crat_31_lr == io_rj_3,
       crat_30_valid & crat_30_lr == io_rj_3,
       crat_29_valid & crat_29_lr == io_rj_3,
       crat_28_valid & crat_28_lr == io_rj_3,
       crat_27_valid & crat_27_lr == io_rj_3,
       crat_26_valid & crat_26_lr == io_rj_3,
       crat_25_valid & crat_25_lr == io_rj_3,
       crat_24_valid & crat_24_lr == io_rj_3,
       crat_23_valid & crat_23_lr == io_rj_3,
       crat_22_valid & crat_22_lr == io_rj_3,
       crat_21_valid & crat_21_lr == io_rj_3,
       crat_20_valid & crat_20_lr == io_rj_3,
       crat_19_valid & crat_19_lr == io_rj_3,
       crat_18_valid & crat_18_lr == io_rj_3,
       crat_17_valid & crat_17_lr == io_rj_3,
       crat_16_valid & crat_16_lr == io_rj_3,
       crat_15_valid & crat_15_lr == io_rj_3,
       crat_14_valid & crat_14_lr == io_rj_3,
       crat_13_valid & crat_13_lr == io_rj_3,
       crat_12_valid & crat_12_lr == io_rj_3,
       crat_11_valid & crat_11_lr == io_rj_3,
       crat_10_valid & crat_10_lr == io_rj_3,
       crat_9_valid & crat_9_lr == io_rj_3,
       crat_8_valid & crat_8_lr == io_rj_3,
       crat_7_valid & crat_7_lr == io_rj_3,
       crat_6_valid & crat_6_lr == io_rj_3,
       crat_5_valid & crat_5_lr == io_rj_3,
       crat_4_valid & crat_4_lr == io_rj_3,
       crat_3_valid & crat_3_lr == io_rj_3,
       crat_2_valid & crat_2_lr == io_rj_3,
       crat_1_valid & crat_1_lr == io_rj_3};
  wire [14:0] _io_prj_3_T_1075 = _io_prj_3_T_1073[30:16] | _io_prj_3_T_1073[14:0];
  wire [6:0]  _io_prj_3_T_1077 = _io_prj_3_T_1075[14:8] | _io_prj_3_T_1075[6:0];
  wire [2:0]  _io_prj_3_T_1079 = _io_prj_3_T_1077[6:4] | _io_prj_3_T_1077[2:0];
  wire [30:0] _io_prk_3_T_1073 =
    {rk_hit_oh_3_63,
     rk_hit_oh_3_62,
     rk_hit_oh_3_61,
     rk_hit_oh_3_60,
     rk_hit_oh_3_59,
     rk_hit_oh_3_58,
     rk_hit_oh_3_57,
     rk_hit_oh_3_56,
     rk_hit_oh_3_55,
     rk_hit_oh_3_54,
     rk_hit_oh_3_53,
     rk_hit_oh_3_52,
     rk_hit_oh_3_51,
     rk_hit_oh_3_50,
     rk_hit_oh_3_49,
     rk_hit_oh_3_48,
     rk_hit_oh_3_47,
     rk_hit_oh_3_46,
     rk_hit_oh_3_45,
     rk_hit_oh_3_44,
     rk_hit_oh_3_43,
     rk_hit_oh_3_42,
     rk_hit_oh_3_41,
     rk_hit_oh_3_40,
     rk_hit_oh_3_39,
     rk_hit_oh_3_38,
     rk_hit_oh_3_37,
     rk_hit_oh_3_36,
     rk_hit_oh_3_35,
     rk_hit_oh_3_34,
     rk_hit_oh_3_33}
    | {crat_31_valid & crat_31_lr == io_rk_3,
       crat_30_valid & crat_30_lr == io_rk_3,
       crat_29_valid & crat_29_lr == io_rk_3,
       crat_28_valid & crat_28_lr == io_rk_3,
       crat_27_valid & crat_27_lr == io_rk_3,
       crat_26_valid & crat_26_lr == io_rk_3,
       crat_25_valid & crat_25_lr == io_rk_3,
       crat_24_valid & crat_24_lr == io_rk_3,
       crat_23_valid & crat_23_lr == io_rk_3,
       crat_22_valid & crat_22_lr == io_rk_3,
       crat_21_valid & crat_21_lr == io_rk_3,
       crat_20_valid & crat_20_lr == io_rk_3,
       crat_19_valid & crat_19_lr == io_rk_3,
       crat_18_valid & crat_18_lr == io_rk_3,
       crat_17_valid & crat_17_lr == io_rk_3,
       crat_16_valid & crat_16_lr == io_rk_3,
       crat_15_valid & crat_15_lr == io_rk_3,
       crat_14_valid & crat_14_lr == io_rk_3,
       crat_13_valid & crat_13_lr == io_rk_3,
       crat_12_valid & crat_12_lr == io_rk_3,
       crat_11_valid & crat_11_lr == io_rk_3,
       crat_10_valid & crat_10_lr == io_rk_3,
       crat_9_valid & crat_9_lr == io_rk_3,
       crat_8_valid & crat_8_lr == io_rk_3,
       crat_7_valid & crat_7_lr == io_rk_3,
       crat_6_valid & crat_6_lr == io_rk_3,
       crat_5_valid & crat_5_lr == io_rk_3,
       crat_4_valid & crat_4_lr == io_rk_3,
       crat_3_valid & crat_3_lr == io_rk_3,
       crat_2_valid & crat_2_lr == io_rk_3,
       crat_1_valid & crat_1_lr == io_rk_3};
  wire [14:0] _io_prk_3_T_1075 = _io_prk_3_T_1073[30:16] | _io_prk_3_T_1073[14:0];
  wire [6:0]  _io_prk_3_T_1077 = _io_prk_3_T_1075[14:8] | _io_prk_3_T_1075[6:0];
  wire [2:0]  _io_prk_3_T_1079 = _io_prk_3_T_1077[6:4] | _io_prk_3_T_1077[2:0];
  wire [30:0] _io_pprd_3_T_1073 =
    {rd_hit_oh_3_63,
     rd_hit_oh_3_62,
     rd_hit_oh_3_61,
     rd_hit_oh_3_60,
     rd_hit_oh_3_59,
     rd_hit_oh_3_58,
     rd_hit_oh_3_57,
     rd_hit_oh_3_56,
     rd_hit_oh_3_55,
     rd_hit_oh_3_54,
     rd_hit_oh_3_53,
     rd_hit_oh_3_52,
     rd_hit_oh_3_51,
     rd_hit_oh_3_50,
     rd_hit_oh_3_49,
     rd_hit_oh_3_48,
     rd_hit_oh_3_47,
     rd_hit_oh_3_46,
     rd_hit_oh_3_45,
     rd_hit_oh_3_44,
     rd_hit_oh_3_43,
     rd_hit_oh_3_42,
     rd_hit_oh_3_41,
     rd_hit_oh_3_40,
     rd_hit_oh_3_39,
     rd_hit_oh_3_38,
     rd_hit_oh_3_37,
     rd_hit_oh_3_36,
     rd_hit_oh_3_35,
     rd_hit_oh_3_34,
     rd_hit_oh_3_33}
    | {crat_31_valid & crat_31_lr == io_rd_3,
       crat_30_valid & crat_30_lr == io_rd_3,
       crat_29_valid & crat_29_lr == io_rd_3,
       crat_28_valid & crat_28_lr == io_rd_3,
       crat_27_valid & crat_27_lr == io_rd_3,
       crat_26_valid & crat_26_lr == io_rd_3,
       crat_25_valid & crat_25_lr == io_rd_3,
       crat_24_valid & crat_24_lr == io_rd_3,
       crat_23_valid & crat_23_lr == io_rd_3,
       crat_22_valid & crat_22_lr == io_rd_3,
       crat_21_valid & crat_21_lr == io_rd_3,
       crat_20_valid & crat_20_lr == io_rd_3,
       crat_19_valid & crat_19_lr == io_rd_3,
       crat_18_valid & crat_18_lr == io_rd_3,
       crat_17_valid & crat_17_lr == io_rd_3,
       crat_16_valid & crat_16_lr == io_rd_3,
       crat_15_valid & crat_15_lr == io_rd_3,
       crat_14_valid & crat_14_lr == io_rd_3,
       crat_13_valid & crat_13_lr == io_rd_3,
       crat_12_valid & crat_12_lr == io_rd_3,
       crat_11_valid & crat_11_lr == io_rd_3,
       crat_10_valid & crat_10_lr == io_rd_3,
       crat_9_valid & crat_9_lr == io_rd_3,
       crat_8_valid & crat_8_lr == io_rd_3,
       crat_7_valid & crat_7_lr == io_rd_3,
       crat_6_valid & crat_6_lr == io_rd_3,
       crat_5_valid & crat_5_lr == io_rd_3,
       crat_4_valid & crat_4_lr == io_rd_3,
       crat_3_valid & crat_3_lr == io_rd_3,
       crat_2_valid & crat_2_lr == io_rd_3,
       crat_1_valid & crat_1_lr == io_rd_3};
  wire [14:0] _io_pprd_3_T_1075 = _io_pprd_3_T_1073[30:16] | _io_pprd_3_T_1073[14:0];
  wire [6:0]  _io_pprd_3_T_1077 = _io_pprd_3_T_1075[14:8] | _io_pprd_3_T_1075[6:0];
  wire [2:0]  _io_pprd_3_T_1079 = _io_pprd_3_T_1077[6:4] | _io_pprd_3_T_1077[2:0];
  wire [5:0]  _io_pprd_3_output =
    {|{rd_hit_oh_3_63,
       rd_hit_oh_3_62,
       rd_hit_oh_3_61,
       rd_hit_oh_3_60,
       rd_hit_oh_3_59,
       rd_hit_oh_3_58,
       rd_hit_oh_3_57,
       rd_hit_oh_3_56,
       rd_hit_oh_3_55,
       rd_hit_oh_3_54,
       rd_hit_oh_3_53,
       rd_hit_oh_3_52,
       rd_hit_oh_3_51,
       rd_hit_oh_3_50,
       rd_hit_oh_3_49,
       rd_hit_oh_3_48,
       rd_hit_oh_3_47,
       rd_hit_oh_3_46,
       rd_hit_oh_3_45,
       rd_hit_oh_3_44,
       rd_hit_oh_3_43,
       rd_hit_oh_3_42,
       rd_hit_oh_3_41,
       rd_hit_oh_3_40,
       rd_hit_oh_3_39,
       rd_hit_oh_3_38,
       rd_hit_oh_3_37,
       rd_hit_oh_3_36,
       rd_hit_oh_3_35,
       rd_hit_oh_3_34,
       rd_hit_oh_3_33,
       crat_32_valid & crat_32_lr == io_rd_3},
     |(_io_pprd_3_T_1073[30:15]),
     |(_io_pprd_3_T_1075[14:7]),
     |(_io_pprd_3_T_1077[6:3]),
     |(_io_pprd_3_T_1079[2:1]),
     _io_pprd_3_T_1079[2] | _io_pprd_3_T_1079[0]};
  wire        _GEN = ~reset & crat_0_valid;
  wire        _GEN_0 = ~reset & crat_1_valid;
  wire        _GEN_1 = ~reset & crat_2_valid;
  wire        _GEN_2 = ~reset & crat_3_valid;
  wire        _GEN_3 = ~reset & crat_4_valid;
  wire        _GEN_4 = ~reset & crat_5_valid;
  wire        _GEN_5 = ~reset & crat_6_valid;
  wire        _GEN_6 = ~reset & crat_7_valid;
  wire        _GEN_7 = ~reset & crat_8_valid;
  wire        _GEN_8 = ~reset & crat_9_valid;
  wire        _GEN_9 = ~reset & crat_10_valid;
  wire        _GEN_10 = ~reset & crat_11_valid;
  wire        _GEN_11 = ~reset & crat_12_valid;
  wire        _GEN_12 = ~reset & crat_13_valid;
  wire        _GEN_13 = ~reset & crat_14_valid;
  wire        _GEN_14 = ~reset & crat_15_valid;
  wire        _GEN_15 = ~reset & crat_16_valid;
  wire        _GEN_16 = ~reset & crat_17_valid;
  wire        _GEN_17 = ~reset & crat_18_valid;
  wire        _GEN_18 = ~reset & crat_19_valid;
  wire        _GEN_19 = ~reset & crat_20_valid;
  wire        _GEN_20 = ~reset & crat_21_valid;
  wire        _GEN_21 = ~reset & crat_22_valid;
  wire        _GEN_22 = ~reset & crat_23_valid;
  wire        _GEN_23 = ~reset & crat_24_valid;
  wire        _GEN_24 = ~reset & crat_25_valid;
  wire        _GEN_25 = ~reset & crat_26_valid;
  wire        _GEN_26 = ~reset & crat_27_valid;
  wire        _GEN_27 = ~reset & crat_28_valid;
  wire        _GEN_28 = ~reset & crat_29_valid;
  wire        _GEN_29 = ~reset & crat_30_valid;
  wire        _GEN_30 = ~reset & crat_31_valid;
  wire        _GEN_31 = ~reset & crat_32_valid;
  wire        _GEN_32 = ~reset & crat_33_valid;
  wire        _GEN_33 = ~reset & crat_34_valid;
  wire        _GEN_34 = ~reset & crat_35_valid;
  wire        _GEN_35 = ~reset & crat_36_valid;
  wire        _GEN_36 = ~reset & crat_37_valid;
  wire        _GEN_37 = ~reset & crat_38_valid;
  wire        _GEN_38 = ~reset & crat_39_valid;
  wire        _GEN_39 = ~reset & crat_40_valid;
  wire        _GEN_40 = ~reset & crat_41_valid;
  wire        _GEN_41 = ~reset & crat_42_valid;
  wire        _GEN_42 = ~reset & crat_43_valid;
  wire        _GEN_43 = ~reset & crat_44_valid;
  wire        _GEN_44 = ~reset & crat_45_valid;
  wire        _GEN_45 = ~reset & crat_46_valid;
  wire        _GEN_46 = ~reset & crat_47_valid;
  wire        _GEN_47 = ~reset & crat_48_valid;
  wire        _GEN_48 = ~reset & crat_49_valid;
  wire        _GEN_49 = ~reset & crat_50_valid;
  wire        _GEN_50 = ~reset & crat_51_valid;
  wire        _GEN_51 = ~reset & crat_52_valid;
  wire        _GEN_52 = ~reset & crat_53_valid;
  wire        _GEN_53 = ~reset & crat_54_valid;
  wire        _GEN_54 = ~reset & crat_55_valid;
  wire        _GEN_55 = ~reset & crat_56_valid;
  wire        _GEN_56 = ~reset & crat_57_valid;
  wire        _GEN_57 = ~reset & crat_58_valid;
  wire        _GEN_58 = ~reset & crat_59_valid;
  wire        _GEN_59 = ~reset & crat_60_valid;
  wire        _GEN_60 = ~reset & crat_61_valid;
  wire        _GEN_61 = ~reset & crat_62_valid;
  wire        _GEN_62 = ~reset & crat_63_valid;
  wire        _GEN_63 = io_alloc_preg_0 == 6'h0;
  wire        _GEN_64 = io_alloc_preg_0 == 6'h1;
  wire        _GEN_65 = io_alloc_preg_0 == 6'h2;
  wire        _GEN_66 = io_alloc_preg_0 == 6'h3;
  wire        _GEN_67 = io_alloc_preg_0 == 6'h4;
  wire        _GEN_68 = io_alloc_preg_0 == 6'h5;
  wire        _GEN_69 = io_alloc_preg_0 == 6'h6;
  wire        _GEN_70 = io_alloc_preg_0 == 6'h7;
  wire        _GEN_71 = io_alloc_preg_0 == 6'h8;
  wire        _GEN_72 = io_alloc_preg_0 == 6'h9;
  wire        _GEN_73 = io_alloc_preg_0 == 6'hA;
  wire        _GEN_74 = io_alloc_preg_0 == 6'hB;
  wire        _GEN_75 = io_alloc_preg_0 == 6'hC;
  wire        _GEN_76 = io_alloc_preg_0 == 6'hD;
  wire        _GEN_77 = io_alloc_preg_0 == 6'hE;
  wire        _GEN_78 = io_alloc_preg_0 == 6'hF;
  wire        _GEN_79 = io_alloc_preg_0 == 6'h10;
  wire        _GEN_80 = io_alloc_preg_0 == 6'h11;
  wire        _GEN_81 = io_alloc_preg_0 == 6'h12;
  wire        _GEN_82 = io_alloc_preg_0 == 6'h13;
  wire        _GEN_83 = io_alloc_preg_0 == 6'h14;
  wire        _GEN_84 = io_alloc_preg_0 == 6'h15;
  wire        _GEN_85 = io_alloc_preg_0 == 6'h16;
  wire        _GEN_86 = io_alloc_preg_0 == 6'h17;
  wire        _GEN_87 = io_alloc_preg_0 == 6'h18;
  wire        _GEN_88 = io_alloc_preg_0 == 6'h19;
  wire        _GEN_89 = io_alloc_preg_0 == 6'h1A;
  wire        _GEN_90 = io_alloc_preg_0 == 6'h1B;
  wire        _GEN_91 = io_alloc_preg_0 == 6'h1C;
  wire        _GEN_92 = io_alloc_preg_0 == 6'h1D;
  wire        _GEN_93 = io_alloc_preg_0 == 6'h1E;
  wire        _GEN_94 = io_alloc_preg_0 == 6'h1F;
  wire        _GEN_95 = io_alloc_preg_0 == 6'h20;
  wire        _GEN_96 = io_alloc_preg_0 == 6'h21;
  wire        _GEN_97 = io_alloc_preg_0 == 6'h22;
  wire        _GEN_98 = io_alloc_preg_0 == 6'h23;
  wire        _GEN_99 = io_alloc_preg_0 == 6'h24;
  wire        _GEN_100 = io_alloc_preg_0 == 6'h25;
  wire        _GEN_101 = io_alloc_preg_0 == 6'h26;
  wire        _GEN_102 = io_alloc_preg_0 == 6'h27;
  wire        _GEN_103 = io_alloc_preg_0 == 6'h28;
  wire        _GEN_104 = io_alloc_preg_0 == 6'h29;
  wire        _GEN_105 = io_alloc_preg_0 == 6'h2A;
  wire        _GEN_106 = io_alloc_preg_0 == 6'h2B;
  wire        _GEN_107 = io_alloc_preg_0 == 6'h2C;
  wire        _GEN_108 = io_alloc_preg_0 == 6'h2D;
  wire        _GEN_109 = io_alloc_preg_0 == 6'h2E;
  wire        _GEN_110 = io_alloc_preg_0 == 6'h2F;
  wire        _GEN_111 = io_alloc_preg_0 == 6'h30;
  wire        _GEN_112 = io_alloc_preg_0 == 6'h31;
  wire        _GEN_113 = io_alloc_preg_0 == 6'h32;
  wire        _GEN_114 = io_alloc_preg_0 == 6'h33;
  wire        _GEN_115 = io_alloc_preg_0 == 6'h34;
  wire        _GEN_116 = io_alloc_preg_0 == 6'h35;
  wire        _GEN_117 = io_alloc_preg_0 == 6'h36;
  wire        _GEN_118 = io_alloc_preg_0 == 6'h37;
  wire        _GEN_119 = io_alloc_preg_0 == 6'h38;
  wire        _GEN_120 = io_alloc_preg_0 == 6'h39;
  wire        _GEN_121 = io_alloc_preg_0 == 6'h3A;
  wire        _GEN_122 = io_alloc_preg_0 == 6'h3B;
  wire        _GEN_123 = io_alloc_preg_0 == 6'h3C;
  wire        _GEN_124 = io_alloc_preg_0 == 6'h3D;
  wire        _GEN_125 = io_alloc_preg_0 == 6'h3E;
  wire        _GEN_126 = (|_io_pprd_0_output) & (_GEN_63 | _GEN);
  wire        _GEN_127 = io_rd_valid_0 ? _GEN_126 : _GEN;
  wire        _GEN_128 = _io_pprd_0_output != 6'h1 & (_GEN_64 | _GEN_0);
  wire        _GEN_129 = io_rd_valid_0 ? _GEN_128 : _GEN_0;
  wire        _GEN_130 = _io_pprd_0_output != 6'h2 & (_GEN_65 | _GEN_1);
  wire        _GEN_131 = io_rd_valid_0 ? _GEN_130 : _GEN_1;
  wire        _GEN_132 = _io_pprd_0_output != 6'h3 & (_GEN_66 | _GEN_2);
  wire        _GEN_133 = io_rd_valid_0 ? _GEN_132 : _GEN_2;
  wire        _GEN_134 = _io_pprd_0_output != 6'h4 & (_GEN_67 | _GEN_3);
  wire        _GEN_135 = io_rd_valid_0 ? _GEN_134 : _GEN_3;
  wire        _GEN_136 = _io_pprd_0_output != 6'h5 & (_GEN_68 | _GEN_4);
  wire        _GEN_137 = io_rd_valid_0 ? _GEN_136 : _GEN_4;
  wire        _GEN_138 = _io_pprd_0_output != 6'h6 & (_GEN_69 | _GEN_5);
  wire        _GEN_139 = io_rd_valid_0 ? _GEN_138 : _GEN_5;
  wire        _GEN_140 = _io_pprd_0_output != 6'h7 & (_GEN_70 | _GEN_6);
  wire        _GEN_141 = io_rd_valid_0 ? _GEN_140 : _GEN_6;
  wire        _GEN_142 = _io_pprd_0_output != 6'h8 & (_GEN_71 | _GEN_7);
  wire        _GEN_143 = io_rd_valid_0 ? _GEN_142 : _GEN_7;
  wire        _GEN_144 = _io_pprd_0_output != 6'h9 & (_GEN_72 | _GEN_8);
  wire        _GEN_145 = io_rd_valid_0 ? _GEN_144 : _GEN_8;
  wire        _GEN_146 = _io_pprd_0_output != 6'hA & (_GEN_73 | _GEN_9);
  wire        _GEN_147 = io_rd_valid_0 ? _GEN_146 : _GEN_9;
  wire        _GEN_148 = _io_pprd_0_output != 6'hB & (_GEN_74 | _GEN_10);
  wire        _GEN_149 = io_rd_valid_0 ? _GEN_148 : _GEN_10;
  wire        _GEN_150 = _io_pprd_0_output != 6'hC & (_GEN_75 | _GEN_11);
  wire        _GEN_151 = io_rd_valid_0 ? _GEN_150 : _GEN_11;
  wire        _GEN_152 = _io_pprd_0_output != 6'hD & (_GEN_76 | _GEN_12);
  wire        _GEN_153 = io_rd_valid_0 ? _GEN_152 : _GEN_12;
  wire        _GEN_154 = _io_pprd_0_output != 6'hE & (_GEN_77 | _GEN_13);
  wire        _GEN_155 = io_rd_valid_0 ? _GEN_154 : _GEN_13;
  wire        _GEN_156 = _io_pprd_0_output != 6'hF & (_GEN_78 | _GEN_14);
  wire        _GEN_157 = io_rd_valid_0 ? _GEN_156 : _GEN_14;
  wire        _GEN_158 = _io_pprd_0_output != 6'h10 & (_GEN_79 | _GEN_15);
  wire        _GEN_159 = io_rd_valid_0 ? _GEN_158 : _GEN_15;
  wire        _GEN_160 = _io_pprd_0_output != 6'h11 & (_GEN_80 | _GEN_16);
  wire        _GEN_161 = io_rd_valid_0 ? _GEN_160 : _GEN_16;
  wire        _GEN_162 = _io_pprd_0_output != 6'h12 & (_GEN_81 | _GEN_17);
  wire        _GEN_163 = io_rd_valid_0 ? _GEN_162 : _GEN_17;
  wire        _GEN_164 = _io_pprd_0_output != 6'h13 & (_GEN_82 | _GEN_18);
  wire        _GEN_165 = io_rd_valid_0 ? _GEN_164 : _GEN_18;
  wire        _GEN_166 = _io_pprd_0_output != 6'h14 & (_GEN_83 | _GEN_19);
  wire        _GEN_167 = io_rd_valid_0 ? _GEN_166 : _GEN_19;
  wire        _GEN_168 = _io_pprd_0_output != 6'h15 & (_GEN_84 | _GEN_20);
  wire        _GEN_169 = io_rd_valid_0 ? _GEN_168 : _GEN_20;
  wire        _GEN_170 = _io_pprd_0_output != 6'h16 & (_GEN_85 | _GEN_21);
  wire        _GEN_171 = io_rd_valid_0 ? _GEN_170 : _GEN_21;
  wire        _GEN_172 = _io_pprd_0_output != 6'h17 & (_GEN_86 | _GEN_22);
  wire        _GEN_173 = io_rd_valid_0 ? _GEN_172 : _GEN_22;
  wire        _GEN_174 = _io_pprd_0_output != 6'h18 & (_GEN_87 | _GEN_23);
  wire        _GEN_175 = io_rd_valid_0 ? _GEN_174 : _GEN_23;
  wire        _GEN_176 = _io_pprd_0_output != 6'h19 & (_GEN_88 | _GEN_24);
  wire        _GEN_177 = io_rd_valid_0 ? _GEN_176 : _GEN_24;
  wire        _GEN_178 = _io_pprd_0_output != 6'h1A & (_GEN_89 | _GEN_25);
  wire        _GEN_179 = io_rd_valid_0 ? _GEN_178 : _GEN_25;
  wire        _GEN_180 = _io_pprd_0_output != 6'h1B & (_GEN_90 | _GEN_26);
  wire        _GEN_181 = io_rd_valid_0 ? _GEN_180 : _GEN_26;
  wire        _GEN_182 = _io_pprd_0_output != 6'h1C & (_GEN_91 | _GEN_27);
  wire        _GEN_183 = io_rd_valid_0 ? _GEN_182 : _GEN_27;
  wire        _GEN_184 = _io_pprd_0_output != 6'h1D & (_GEN_92 | _GEN_28);
  wire        _GEN_185 = io_rd_valid_0 ? _GEN_184 : _GEN_28;
  wire        _GEN_186 = _io_pprd_0_output != 6'h1E & (_GEN_93 | _GEN_29);
  wire        _GEN_187 = io_rd_valid_0 ? _GEN_186 : _GEN_29;
  wire        _GEN_188 = _io_pprd_0_output != 6'h1F & (_GEN_94 | _GEN_30);
  wire        _GEN_189 = io_rd_valid_0 ? _GEN_188 : _GEN_30;
  wire        _GEN_190 = _io_pprd_0_output != 6'h20 & (_GEN_95 | _GEN_31);
  wire        _GEN_191 = io_rd_valid_0 ? _GEN_190 : _GEN_31;
  wire        _GEN_192 = _io_pprd_0_output != 6'h21 & (_GEN_96 | _GEN_32);
  wire        _GEN_193 = io_rd_valid_0 ? _GEN_192 : _GEN_32;
  wire        _GEN_194 = _io_pprd_0_output != 6'h22 & (_GEN_97 | _GEN_33);
  wire        _GEN_195 = io_rd_valid_0 ? _GEN_194 : _GEN_33;
  wire        _GEN_196 = _io_pprd_0_output != 6'h23 & (_GEN_98 | _GEN_34);
  wire        _GEN_197 = io_rd_valid_0 ? _GEN_196 : _GEN_34;
  wire        _GEN_198 = _io_pprd_0_output != 6'h24 & (_GEN_99 | _GEN_35);
  wire        _GEN_199 = io_rd_valid_0 ? _GEN_198 : _GEN_35;
  wire        _GEN_200 = _io_pprd_0_output != 6'h25 & (_GEN_100 | _GEN_36);
  wire        _GEN_201 = io_rd_valid_0 ? _GEN_200 : _GEN_36;
  wire        _GEN_202 = _io_pprd_0_output != 6'h26 & (_GEN_101 | _GEN_37);
  wire        _GEN_203 = io_rd_valid_0 ? _GEN_202 : _GEN_37;
  wire        _GEN_204 = _io_pprd_0_output != 6'h27 & (_GEN_102 | _GEN_38);
  wire        _GEN_205 = io_rd_valid_0 ? _GEN_204 : _GEN_38;
  wire        _GEN_206 = _io_pprd_0_output != 6'h28 & (_GEN_103 | _GEN_39);
  wire        _GEN_207 = io_rd_valid_0 ? _GEN_206 : _GEN_39;
  wire        _GEN_208 = _io_pprd_0_output != 6'h29 & (_GEN_104 | _GEN_40);
  wire        _GEN_209 = io_rd_valid_0 ? _GEN_208 : _GEN_40;
  wire        _GEN_210 = _io_pprd_0_output != 6'h2A & (_GEN_105 | _GEN_41);
  wire        _GEN_211 = io_rd_valid_0 ? _GEN_210 : _GEN_41;
  wire        _GEN_212 = _io_pprd_0_output != 6'h2B & (_GEN_106 | _GEN_42);
  wire        _GEN_213 = io_rd_valid_0 ? _GEN_212 : _GEN_42;
  wire        _GEN_214 = _io_pprd_0_output != 6'h2C & (_GEN_107 | _GEN_43);
  wire        _GEN_215 = io_rd_valid_0 ? _GEN_214 : _GEN_43;
  wire        _GEN_216 = _io_pprd_0_output != 6'h2D & (_GEN_108 | _GEN_44);
  wire        _GEN_217 = io_rd_valid_0 ? _GEN_216 : _GEN_44;
  wire        _GEN_218 = _io_pprd_0_output != 6'h2E & (_GEN_109 | _GEN_45);
  wire        _GEN_219 = io_rd_valid_0 ? _GEN_218 : _GEN_45;
  wire        _GEN_220 = _io_pprd_0_output != 6'h2F & (_GEN_110 | _GEN_46);
  wire        _GEN_221 = io_rd_valid_0 ? _GEN_220 : _GEN_46;
  wire        _GEN_222 = _io_pprd_0_output != 6'h30 & (_GEN_111 | _GEN_47);
  wire        _GEN_223 = io_rd_valid_0 ? _GEN_222 : _GEN_47;
  wire        _GEN_224 = _io_pprd_0_output != 6'h31 & (_GEN_112 | _GEN_48);
  wire        _GEN_225 = io_rd_valid_0 ? _GEN_224 : _GEN_48;
  wire        _GEN_226 = _io_pprd_0_output != 6'h32 & (_GEN_113 | _GEN_49);
  wire        _GEN_227 = io_rd_valid_0 ? _GEN_226 : _GEN_49;
  wire        _GEN_228 = _io_pprd_0_output != 6'h33 & (_GEN_114 | _GEN_50);
  wire        _GEN_229 = io_rd_valid_0 ? _GEN_228 : _GEN_50;
  wire        _GEN_230 = _io_pprd_0_output != 6'h34 & (_GEN_115 | _GEN_51);
  wire        _GEN_231 = io_rd_valid_0 ? _GEN_230 : _GEN_51;
  wire        _GEN_232 = _io_pprd_0_output != 6'h35 & (_GEN_116 | _GEN_52);
  wire        _GEN_233 = io_rd_valid_0 ? _GEN_232 : _GEN_52;
  wire        _GEN_234 = _io_pprd_0_output != 6'h36 & (_GEN_117 | _GEN_53);
  wire        _GEN_235 = io_rd_valid_0 ? _GEN_234 : _GEN_53;
  wire        _GEN_236 = _io_pprd_0_output != 6'h37 & (_GEN_118 | _GEN_54);
  wire        _GEN_237 = io_rd_valid_0 ? _GEN_236 : _GEN_54;
  wire        _GEN_238 = _io_pprd_0_output != 6'h38 & (_GEN_119 | _GEN_55);
  wire        _GEN_239 = io_rd_valid_0 ? _GEN_238 : _GEN_55;
  wire        _GEN_240 = _io_pprd_0_output != 6'h39 & (_GEN_120 | _GEN_56);
  wire        _GEN_241 = io_rd_valid_0 ? _GEN_240 : _GEN_56;
  wire        _GEN_242 = _io_pprd_0_output != 6'h3A & (_GEN_121 | _GEN_57);
  wire        _GEN_243 = io_rd_valid_0 ? _GEN_242 : _GEN_57;
  wire        _GEN_244 = _io_pprd_0_output != 6'h3B & (_GEN_122 | _GEN_58);
  wire        _GEN_245 = io_rd_valid_0 ? _GEN_244 : _GEN_58;
  wire        _GEN_246 = _io_pprd_0_output != 6'h3C & (_GEN_123 | _GEN_59);
  wire        _GEN_247 = io_rd_valid_0 ? _GEN_246 : _GEN_59;
  wire        _GEN_248 = _io_pprd_0_output != 6'h3D & (_GEN_124 | _GEN_60);
  wire        _GEN_249 = io_rd_valid_0 ? _GEN_248 : _GEN_60;
  wire        _GEN_250 = _io_pprd_0_output != 6'h3E & (_GEN_125 | _GEN_61);
  wire        _GEN_251 = io_rd_valid_0 ? _GEN_250 : _GEN_61;
  wire        _GEN_252 = _io_pprd_0_output != 6'h3F & ((&io_alloc_preg_0) | _GEN_62);
  wire        _GEN_253 = io_rd_valid_0 ? _GEN_252 : _GEN_62;
  wire        _GEN_254 = io_alloc_preg_1 == 6'h0;
  wire        _GEN_255 = io_alloc_preg_1 == 6'h1;
  wire        _GEN_256 = io_alloc_preg_1 == 6'h2;
  wire        _GEN_257 = io_alloc_preg_1 == 6'h3;
  wire        _GEN_258 = io_alloc_preg_1 == 6'h4;
  wire        _GEN_259 = io_alloc_preg_1 == 6'h5;
  wire        _GEN_260 = io_alloc_preg_1 == 6'h6;
  wire        _GEN_261 = io_alloc_preg_1 == 6'h7;
  wire        _GEN_262 = io_alloc_preg_1 == 6'h8;
  wire        _GEN_263 = io_alloc_preg_1 == 6'h9;
  wire        _GEN_264 = io_alloc_preg_1 == 6'hA;
  wire        _GEN_265 = io_alloc_preg_1 == 6'hB;
  wire        _GEN_266 = io_alloc_preg_1 == 6'hC;
  wire        _GEN_267 = io_alloc_preg_1 == 6'hD;
  wire        _GEN_268 = io_alloc_preg_1 == 6'hE;
  wire        _GEN_269 = io_alloc_preg_1 == 6'hF;
  wire        _GEN_270 = io_alloc_preg_1 == 6'h10;
  wire        _GEN_271 = io_alloc_preg_1 == 6'h11;
  wire        _GEN_272 = io_alloc_preg_1 == 6'h12;
  wire        _GEN_273 = io_alloc_preg_1 == 6'h13;
  wire        _GEN_274 = io_alloc_preg_1 == 6'h14;
  wire        _GEN_275 = io_alloc_preg_1 == 6'h15;
  wire        _GEN_276 = io_alloc_preg_1 == 6'h16;
  wire        _GEN_277 = io_alloc_preg_1 == 6'h17;
  wire        _GEN_278 = io_alloc_preg_1 == 6'h18;
  wire        _GEN_279 = io_alloc_preg_1 == 6'h19;
  wire        _GEN_280 = io_alloc_preg_1 == 6'h1A;
  wire        _GEN_281 = io_alloc_preg_1 == 6'h1B;
  wire        _GEN_282 = io_alloc_preg_1 == 6'h1C;
  wire        _GEN_283 = io_alloc_preg_1 == 6'h1D;
  wire        _GEN_284 = io_alloc_preg_1 == 6'h1E;
  wire        _GEN_285 = io_alloc_preg_1 == 6'h1F;
  wire        _GEN_286 = io_alloc_preg_1 == 6'h20;
  wire        _GEN_287 = io_alloc_preg_1 == 6'h21;
  wire        _GEN_288 = io_alloc_preg_1 == 6'h22;
  wire        _GEN_289 = io_alloc_preg_1 == 6'h23;
  wire        _GEN_290 = io_alloc_preg_1 == 6'h24;
  wire        _GEN_291 = io_alloc_preg_1 == 6'h25;
  wire        _GEN_292 = io_alloc_preg_1 == 6'h26;
  wire        _GEN_293 = io_alloc_preg_1 == 6'h27;
  wire        _GEN_294 = io_alloc_preg_1 == 6'h28;
  wire        _GEN_295 = io_alloc_preg_1 == 6'h29;
  wire        _GEN_296 = io_alloc_preg_1 == 6'h2A;
  wire        _GEN_297 = io_alloc_preg_1 == 6'h2B;
  wire        _GEN_298 = io_alloc_preg_1 == 6'h2C;
  wire        _GEN_299 = io_alloc_preg_1 == 6'h2D;
  wire        _GEN_300 = io_alloc_preg_1 == 6'h2E;
  wire        _GEN_301 = io_alloc_preg_1 == 6'h2F;
  wire        _GEN_302 = io_alloc_preg_1 == 6'h30;
  wire        _GEN_303 = io_alloc_preg_1 == 6'h31;
  wire        _GEN_304 = io_alloc_preg_1 == 6'h32;
  wire        _GEN_305 = io_alloc_preg_1 == 6'h33;
  wire        _GEN_306 = io_alloc_preg_1 == 6'h34;
  wire        _GEN_307 = io_alloc_preg_1 == 6'h35;
  wire        _GEN_308 = io_alloc_preg_1 == 6'h36;
  wire        _GEN_309 = io_alloc_preg_1 == 6'h37;
  wire        _GEN_310 = io_alloc_preg_1 == 6'h38;
  wire        _GEN_311 = io_alloc_preg_1 == 6'h39;
  wire        _GEN_312 = io_alloc_preg_1 == 6'h3A;
  wire        _GEN_313 = io_alloc_preg_1 == 6'h3B;
  wire        _GEN_314 = io_alloc_preg_1 == 6'h3C;
  wire        _GEN_315 = io_alloc_preg_1 == 6'h3D;
  wire        _GEN_316 = io_alloc_preg_1 == 6'h3E;
  wire        _GEN_317 = (|_io_pprd_1_output) & (_GEN_254 | _GEN_127);
  wire        _GEN_318 = io_rd_valid_1 ? _GEN_317 : _GEN_127;
  wire        _GEN_319 = _io_pprd_1_output != 6'h1 & (_GEN_255 | _GEN_129);
  wire        _GEN_320 = io_rd_valid_1 ? _GEN_319 : _GEN_129;
  wire        _GEN_321 = _io_pprd_1_output != 6'h2 & (_GEN_256 | _GEN_131);
  wire        _GEN_322 = io_rd_valid_1 ? _GEN_321 : _GEN_131;
  wire        _GEN_323 = _io_pprd_1_output != 6'h3 & (_GEN_257 | _GEN_133);
  wire        _GEN_324 = io_rd_valid_1 ? _GEN_323 : _GEN_133;
  wire        _GEN_325 = _io_pprd_1_output != 6'h4 & (_GEN_258 | _GEN_135);
  wire        _GEN_326 = io_rd_valid_1 ? _GEN_325 : _GEN_135;
  wire        _GEN_327 = _io_pprd_1_output != 6'h5 & (_GEN_259 | _GEN_137);
  wire        _GEN_328 = io_rd_valid_1 ? _GEN_327 : _GEN_137;
  wire        _GEN_329 = _io_pprd_1_output != 6'h6 & (_GEN_260 | _GEN_139);
  wire        _GEN_330 = io_rd_valid_1 ? _GEN_329 : _GEN_139;
  wire        _GEN_331 = _io_pprd_1_output != 6'h7 & (_GEN_261 | _GEN_141);
  wire        _GEN_332 = io_rd_valid_1 ? _GEN_331 : _GEN_141;
  wire        _GEN_333 = _io_pprd_1_output != 6'h8 & (_GEN_262 | _GEN_143);
  wire        _GEN_334 = io_rd_valid_1 ? _GEN_333 : _GEN_143;
  wire        _GEN_335 = _io_pprd_1_output != 6'h9 & (_GEN_263 | _GEN_145);
  wire        _GEN_336 = io_rd_valid_1 ? _GEN_335 : _GEN_145;
  wire        _GEN_337 = _io_pprd_1_output != 6'hA & (_GEN_264 | _GEN_147);
  wire        _GEN_338 = io_rd_valid_1 ? _GEN_337 : _GEN_147;
  wire        _GEN_339 = _io_pprd_1_output != 6'hB & (_GEN_265 | _GEN_149);
  wire        _GEN_340 = io_rd_valid_1 ? _GEN_339 : _GEN_149;
  wire        _GEN_341 = _io_pprd_1_output != 6'hC & (_GEN_266 | _GEN_151);
  wire        _GEN_342 = io_rd_valid_1 ? _GEN_341 : _GEN_151;
  wire        _GEN_343 = _io_pprd_1_output != 6'hD & (_GEN_267 | _GEN_153);
  wire        _GEN_344 = io_rd_valid_1 ? _GEN_343 : _GEN_153;
  wire        _GEN_345 = _io_pprd_1_output != 6'hE & (_GEN_268 | _GEN_155);
  wire        _GEN_346 = io_rd_valid_1 ? _GEN_345 : _GEN_155;
  wire        _GEN_347 = _io_pprd_1_output != 6'hF & (_GEN_269 | _GEN_157);
  wire        _GEN_348 = io_rd_valid_1 ? _GEN_347 : _GEN_157;
  wire        _GEN_349 = _io_pprd_1_output != 6'h10 & (_GEN_270 | _GEN_159);
  wire        _GEN_350 = io_rd_valid_1 ? _GEN_349 : _GEN_159;
  wire        _GEN_351 = _io_pprd_1_output != 6'h11 & (_GEN_271 | _GEN_161);
  wire        _GEN_352 = io_rd_valid_1 ? _GEN_351 : _GEN_161;
  wire        _GEN_353 = _io_pprd_1_output != 6'h12 & (_GEN_272 | _GEN_163);
  wire        _GEN_354 = io_rd_valid_1 ? _GEN_353 : _GEN_163;
  wire        _GEN_355 = _io_pprd_1_output != 6'h13 & (_GEN_273 | _GEN_165);
  wire        _GEN_356 = io_rd_valid_1 ? _GEN_355 : _GEN_165;
  wire        _GEN_357 = _io_pprd_1_output != 6'h14 & (_GEN_274 | _GEN_167);
  wire        _GEN_358 = io_rd_valid_1 ? _GEN_357 : _GEN_167;
  wire        _GEN_359 = _io_pprd_1_output != 6'h15 & (_GEN_275 | _GEN_169);
  wire        _GEN_360 = io_rd_valid_1 ? _GEN_359 : _GEN_169;
  wire        _GEN_361 = _io_pprd_1_output != 6'h16 & (_GEN_276 | _GEN_171);
  wire        _GEN_362 = io_rd_valid_1 ? _GEN_361 : _GEN_171;
  wire        _GEN_363 = _io_pprd_1_output != 6'h17 & (_GEN_277 | _GEN_173);
  wire        _GEN_364 = io_rd_valid_1 ? _GEN_363 : _GEN_173;
  wire        _GEN_365 = _io_pprd_1_output != 6'h18 & (_GEN_278 | _GEN_175);
  wire        _GEN_366 = io_rd_valid_1 ? _GEN_365 : _GEN_175;
  wire        _GEN_367 = _io_pprd_1_output != 6'h19 & (_GEN_279 | _GEN_177);
  wire        _GEN_368 = io_rd_valid_1 ? _GEN_367 : _GEN_177;
  wire        _GEN_369 = _io_pprd_1_output != 6'h1A & (_GEN_280 | _GEN_179);
  wire        _GEN_370 = io_rd_valid_1 ? _GEN_369 : _GEN_179;
  wire        _GEN_371 = _io_pprd_1_output != 6'h1B & (_GEN_281 | _GEN_181);
  wire        _GEN_372 = io_rd_valid_1 ? _GEN_371 : _GEN_181;
  wire        _GEN_373 = _io_pprd_1_output != 6'h1C & (_GEN_282 | _GEN_183);
  wire        _GEN_374 = io_rd_valid_1 ? _GEN_373 : _GEN_183;
  wire        _GEN_375 = _io_pprd_1_output != 6'h1D & (_GEN_283 | _GEN_185);
  wire        _GEN_376 = io_rd_valid_1 ? _GEN_375 : _GEN_185;
  wire        _GEN_377 = _io_pprd_1_output != 6'h1E & (_GEN_284 | _GEN_187);
  wire        _GEN_378 = io_rd_valid_1 ? _GEN_377 : _GEN_187;
  wire        _GEN_379 = _io_pprd_1_output != 6'h1F & (_GEN_285 | _GEN_189);
  wire        _GEN_380 = io_rd_valid_1 ? _GEN_379 : _GEN_189;
  wire        _GEN_381 = _io_pprd_1_output != 6'h20 & (_GEN_286 | _GEN_191);
  wire        _GEN_382 = io_rd_valid_1 ? _GEN_381 : _GEN_191;
  wire        _GEN_383 = _io_pprd_1_output != 6'h21 & (_GEN_287 | _GEN_193);
  wire        _GEN_384 = io_rd_valid_1 ? _GEN_383 : _GEN_193;
  wire        _GEN_385 = _io_pprd_1_output != 6'h22 & (_GEN_288 | _GEN_195);
  wire        _GEN_386 = io_rd_valid_1 ? _GEN_385 : _GEN_195;
  wire        _GEN_387 = _io_pprd_1_output != 6'h23 & (_GEN_289 | _GEN_197);
  wire        _GEN_388 = io_rd_valid_1 ? _GEN_387 : _GEN_197;
  wire        _GEN_389 = _io_pprd_1_output != 6'h24 & (_GEN_290 | _GEN_199);
  wire        _GEN_390 = io_rd_valid_1 ? _GEN_389 : _GEN_199;
  wire        _GEN_391 = _io_pprd_1_output != 6'h25 & (_GEN_291 | _GEN_201);
  wire        _GEN_392 = io_rd_valid_1 ? _GEN_391 : _GEN_201;
  wire        _GEN_393 = _io_pprd_1_output != 6'h26 & (_GEN_292 | _GEN_203);
  wire        _GEN_394 = io_rd_valid_1 ? _GEN_393 : _GEN_203;
  wire        _GEN_395 = _io_pprd_1_output != 6'h27 & (_GEN_293 | _GEN_205);
  wire        _GEN_396 = io_rd_valid_1 ? _GEN_395 : _GEN_205;
  wire        _GEN_397 = _io_pprd_1_output != 6'h28 & (_GEN_294 | _GEN_207);
  wire        _GEN_398 = io_rd_valid_1 ? _GEN_397 : _GEN_207;
  wire        _GEN_399 = _io_pprd_1_output != 6'h29 & (_GEN_295 | _GEN_209);
  wire        _GEN_400 = io_rd_valid_1 ? _GEN_399 : _GEN_209;
  wire        _GEN_401 = _io_pprd_1_output != 6'h2A & (_GEN_296 | _GEN_211);
  wire        _GEN_402 = io_rd_valid_1 ? _GEN_401 : _GEN_211;
  wire        _GEN_403 = _io_pprd_1_output != 6'h2B & (_GEN_297 | _GEN_213);
  wire        _GEN_404 = io_rd_valid_1 ? _GEN_403 : _GEN_213;
  wire        _GEN_405 = _io_pprd_1_output != 6'h2C & (_GEN_298 | _GEN_215);
  wire        _GEN_406 = io_rd_valid_1 ? _GEN_405 : _GEN_215;
  wire        _GEN_407 = _io_pprd_1_output != 6'h2D & (_GEN_299 | _GEN_217);
  wire        _GEN_408 = io_rd_valid_1 ? _GEN_407 : _GEN_217;
  wire        _GEN_409 = _io_pprd_1_output != 6'h2E & (_GEN_300 | _GEN_219);
  wire        _GEN_410 = io_rd_valid_1 ? _GEN_409 : _GEN_219;
  wire        _GEN_411 = _io_pprd_1_output != 6'h2F & (_GEN_301 | _GEN_221);
  wire        _GEN_412 = io_rd_valid_1 ? _GEN_411 : _GEN_221;
  wire        _GEN_413 = _io_pprd_1_output != 6'h30 & (_GEN_302 | _GEN_223);
  wire        _GEN_414 = io_rd_valid_1 ? _GEN_413 : _GEN_223;
  wire        _GEN_415 = _io_pprd_1_output != 6'h31 & (_GEN_303 | _GEN_225);
  wire        _GEN_416 = io_rd_valid_1 ? _GEN_415 : _GEN_225;
  wire        _GEN_417 = _io_pprd_1_output != 6'h32 & (_GEN_304 | _GEN_227);
  wire        _GEN_418 = io_rd_valid_1 ? _GEN_417 : _GEN_227;
  wire        _GEN_419 = _io_pprd_1_output != 6'h33 & (_GEN_305 | _GEN_229);
  wire        _GEN_420 = io_rd_valid_1 ? _GEN_419 : _GEN_229;
  wire        _GEN_421 = _io_pprd_1_output != 6'h34 & (_GEN_306 | _GEN_231);
  wire        _GEN_422 = io_rd_valid_1 ? _GEN_421 : _GEN_231;
  wire        _GEN_423 = _io_pprd_1_output != 6'h35 & (_GEN_307 | _GEN_233);
  wire        _GEN_424 = io_rd_valid_1 ? _GEN_423 : _GEN_233;
  wire        _GEN_425 = _io_pprd_1_output != 6'h36 & (_GEN_308 | _GEN_235);
  wire        _GEN_426 = io_rd_valid_1 ? _GEN_425 : _GEN_235;
  wire        _GEN_427 = _io_pprd_1_output != 6'h37 & (_GEN_309 | _GEN_237);
  wire        _GEN_428 = io_rd_valid_1 ? _GEN_427 : _GEN_237;
  wire        _GEN_429 = _io_pprd_1_output != 6'h38 & (_GEN_310 | _GEN_239);
  wire        _GEN_430 = io_rd_valid_1 ? _GEN_429 : _GEN_239;
  wire        _GEN_431 = _io_pprd_1_output != 6'h39 & (_GEN_311 | _GEN_241);
  wire        _GEN_432 = io_rd_valid_1 ? _GEN_431 : _GEN_241;
  wire        _GEN_433 = _io_pprd_1_output != 6'h3A & (_GEN_312 | _GEN_243);
  wire        _GEN_434 = io_rd_valid_1 ? _GEN_433 : _GEN_243;
  wire        _GEN_435 = _io_pprd_1_output != 6'h3B & (_GEN_313 | _GEN_245);
  wire        _GEN_436 = io_rd_valid_1 ? _GEN_435 : _GEN_245;
  wire        _GEN_437 = _io_pprd_1_output != 6'h3C & (_GEN_314 | _GEN_247);
  wire        _GEN_438 = io_rd_valid_1 ? _GEN_437 : _GEN_247;
  wire        _GEN_439 = _io_pprd_1_output != 6'h3D & (_GEN_315 | _GEN_249);
  wire        _GEN_440 = io_rd_valid_1 ? _GEN_439 : _GEN_249;
  wire        _GEN_441 = _io_pprd_1_output != 6'h3E & (_GEN_316 | _GEN_251);
  wire        _GEN_442 = io_rd_valid_1 ? _GEN_441 : _GEN_251;
  wire        _GEN_443 = _io_pprd_1_output != 6'h3F & ((&io_alloc_preg_1) | _GEN_253);
  wire        _GEN_444 = io_rd_valid_1 ? _GEN_443 : _GEN_253;
  wire        _GEN_445 = io_alloc_preg_2 == 6'h0;
  wire        _GEN_446 = io_alloc_preg_2 == 6'h1;
  wire        _GEN_447 = io_alloc_preg_2 == 6'h2;
  wire        _GEN_448 = io_alloc_preg_2 == 6'h3;
  wire        _GEN_449 = io_alloc_preg_2 == 6'h4;
  wire        _GEN_450 = io_alloc_preg_2 == 6'h5;
  wire        _GEN_451 = io_alloc_preg_2 == 6'h6;
  wire        _GEN_452 = io_alloc_preg_2 == 6'h7;
  wire        _GEN_453 = io_alloc_preg_2 == 6'h8;
  wire        _GEN_454 = io_alloc_preg_2 == 6'h9;
  wire        _GEN_455 = io_alloc_preg_2 == 6'hA;
  wire        _GEN_456 = io_alloc_preg_2 == 6'hB;
  wire        _GEN_457 = io_alloc_preg_2 == 6'hC;
  wire        _GEN_458 = io_alloc_preg_2 == 6'hD;
  wire        _GEN_459 = io_alloc_preg_2 == 6'hE;
  wire        _GEN_460 = io_alloc_preg_2 == 6'hF;
  wire        _GEN_461 = io_alloc_preg_2 == 6'h10;
  wire        _GEN_462 = io_alloc_preg_2 == 6'h11;
  wire        _GEN_463 = io_alloc_preg_2 == 6'h12;
  wire        _GEN_464 = io_alloc_preg_2 == 6'h13;
  wire        _GEN_465 = io_alloc_preg_2 == 6'h14;
  wire        _GEN_466 = io_alloc_preg_2 == 6'h15;
  wire        _GEN_467 = io_alloc_preg_2 == 6'h16;
  wire        _GEN_468 = io_alloc_preg_2 == 6'h17;
  wire        _GEN_469 = io_alloc_preg_2 == 6'h18;
  wire        _GEN_470 = io_alloc_preg_2 == 6'h19;
  wire        _GEN_471 = io_alloc_preg_2 == 6'h1A;
  wire        _GEN_472 = io_alloc_preg_2 == 6'h1B;
  wire        _GEN_473 = io_alloc_preg_2 == 6'h1C;
  wire        _GEN_474 = io_alloc_preg_2 == 6'h1D;
  wire        _GEN_475 = io_alloc_preg_2 == 6'h1E;
  wire        _GEN_476 = io_alloc_preg_2 == 6'h1F;
  wire        _GEN_477 = io_alloc_preg_2 == 6'h20;
  wire        _GEN_478 = io_alloc_preg_2 == 6'h21;
  wire        _GEN_479 = io_alloc_preg_2 == 6'h22;
  wire        _GEN_480 = io_alloc_preg_2 == 6'h23;
  wire        _GEN_481 = io_alloc_preg_2 == 6'h24;
  wire        _GEN_482 = io_alloc_preg_2 == 6'h25;
  wire        _GEN_483 = io_alloc_preg_2 == 6'h26;
  wire        _GEN_484 = io_alloc_preg_2 == 6'h27;
  wire        _GEN_485 = io_alloc_preg_2 == 6'h28;
  wire        _GEN_486 = io_alloc_preg_2 == 6'h29;
  wire        _GEN_487 = io_alloc_preg_2 == 6'h2A;
  wire        _GEN_488 = io_alloc_preg_2 == 6'h2B;
  wire        _GEN_489 = io_alloc_preg_2 == 6'h2C;
  wire        _GEN_490 = io_alloc_preg_2 == 6'h2D;
  wire        _GEN_491 = io_alloc_preg_2 == 6'h2E;
  wire        _GEN_492 = io_alloc_preg_2 == 6'h2F;
  wire        _GEN_493 = io_alloc_preg_2 == 6'h30;
  wire        _GEN_494 = io_alloc_preg_2 == 6'h31;
  wire        _GEN_495 = io_alloc_preg_2 == 6'h32;
  wire        _GEN_496 = io_alloc_preg_2 == 6'h33;
  wire        _GEN_497 = io_alloc_preg_2 == 6'h34;
  wire        _GEN_498 = io_alloc_preg_2 == 6'h35;
  wire        _GEN_499 = io_alloc_preg_2 == 6'h36;
  wire        _GEN_500 = io_alloc_preg_2 == 6'h37;
  wire        _GEN_501 = io_alloc_preg_2 == 6'h38;
  wire        _GEN_502 = io_alloc_preg_2 == 6'h39;
  wire        _GEN_503 = io_alloc_preg_2 == 6'h3A;
  wire        _GEN_504 = io_alloc_preg_2 == 6'h3B;
  wire        _GEN_505 = io_alloc_preg_2 == 6'h3C;
  wire        _GEN_506 = io_alloc_preg_2 == 6'h3D;
  wire        _GEN_507 = io_alloc_preg_2 == 6'h3E;
  wire        _GEN_508 = (|_io_pprd_2_output) & (_GEN_445 | _GEN_318);
  wire        _GEN_509 = _io_pprd_2_output != 6'h1 & (_GEN_446 | _GEN_320);
  wire        _GEN_510 = _io_pprd_2_output != 6'h2 & (_GEN_447 | _GEN_322);
  wire        _GEN_511 = _io_pprd_2_output != 6'h3 & (_GEN_448 | _GEN_324);
  wire        _GEN_512 = _io_pprd_2_output != 6'h4 & (_GEN_449 | _GEN_326);
  wire        _GEN_513 = _io_pprd_2_output != 6'h5 & (_GEN_450 | _GEN_328);
  wire        _GEN_514 = _io_pprd_2_output != 6'h6 & (_GEN_451 | _GEN_330);
  wire        _GEN_515 = _io_pprd_2_output != 6'h7 & (_GEN_452 | _GEN_332);
  wire        _GEN_516 = _io_pprd_2_output != 6'h8 & (_GEN_453 | _GEN_334);
  wire        _GEN_517 = _io_pprd_2_output != 6'h9 & (_GEN_454 | _GEN_336);
  wire        _GEN_518 = _io_pprd_2_output != 6'hA & (_GEN_455 | _GEN_338);
  wire        _GEN_519 = _io_pprd_2_output != 6'hB & (_GEN_456 | _GEN_340);
  wire        _GEN_520 = _io_pprd_2_output != 6'hC & (_GEN_457 | _GEN_342);
  wire        _GEN_521 = _io_pprd_2_output != 6'hD & (_GEN_458 | _GEN_344);
  wire        _GEN_522 = _io_pprd_2_output != 6'hE & (_GEN_459 | _GEN_346);
  wire        _GEN_523 = _io_pprd_2_output != 6'hF & (_GEN_460 | _GEN_348);
  wire        _GEN_524 = _io_pprd_2_output != 6'h10 & (_GEN_461 | _GEN_350);
  wire        _GEN_525 = _io_pprd_2_output != 6'h11 & (_GEN_462 | _GEN_352);
  wire        _GEN_526 = _io_pprd_2_output != 6'h12 & (_GEN_463 | _GEN_354);
  wire        _GEN_527 = _io_pprd_2_output != 6'h13 & (_GEN_464 | _GEN_356);
  wire        _GEN_528 = _io_pprd_2_output != 6'h14 & (_GEN_465 | _GEN_358);
  wire        _GEN_529 = _io_pprd_2_output != 6'h15 & (_GEN_466 | _GEN_360);
  wire        _GEN_530 = _io_pprd_2_output != 6'h16 & (_GEN_467 | _GEN_362);
  wire        _GEN_531 = _io_pprd_2_output != 6'h17 & (_GEN_468 | _GEN_364);
  wire        _GEN_532 = _io_pprd_2_output != 6'h18 & (_GEN_469 | _GEN_366);
  wire        _GEN_533 = _io_pprd_2_output != 6'h19 & (_GEN_470 | _GEN_368);
  wire        _GEN_534 = _io_pprd_2_output != 6'h1A & (_GEN_471 | _GEN_370);
  wire        _GEN_535 = _io_pprd_2_output != 6'h1B & (_GEN_472 | _GEN_372);
  wire        _GEN_536 = _io_pprd_2_output != 6'h1C & (_GEN_473 | _GEN_374);
  wire        _GEN_537 = _io_pprd_2_output != 6'h1D & (_GEN_474 | _GEN_376);
  wire        _GEN_538 = _io_pprd_2_output != 6'h1E & (_GEN_475 | _GEN_378);
  wire        _GEN_539 = _io_pprd_2_output != 6'h1F & (_GEN_476 | _GEN_380);
  wire        _GEN_540 = _io_pprd_2_output != 6'h20 & (_GEN_477 | _GEN_382);
  wire        _GEN_541 = _io_pprd_2_output != 6'h21 & (_GEN_478 | _GEN_384);
  wire        _GEN_542 = _io_pprd_2_output != 6'h22 & (_GEN_479 | _GEN_386);
  wire        _GEN_543 = _io_pprd_2_output != 6'h23 & (_GEN_480 | _GEN_388);
  wire        _GEN_544 = _io_pprd_2_output != 6'h24 & (_GEN_481 | _GEN_390);
  wire        _GEN_545 = _io_pprd_2_output != 6'h25 & (_GEN_482 | _GEN_392);
  wire        _GEN_546 = _io_pprd_2_output != 6'h26 & (_GEN_483 | _GEN_394);
  wire        _GEN_547 = _io_pprd_2_output != 6'h27 & (_GEN_484 | _GEN_396);
  wire        _GEN_548 = _io_pprd_2_output != 6'h28 & (_GEN_485 | _GEN_398);
  wire        _GEN_549 = _io_pprd_2_output != 6'h29 & (_GEN_486 | _GEN_400);
  wire        _GEN_550 = _io_pprd_2_output != 6'h2A & (_GEN_487 | _GEN_402);
  wire        _GEN_551 = _io_pprd_2_output != 6'h2B & (_GEN_488 | _GEN_404);
  wire        _GEN_552 = _io_pprd_2_output != 6'h2C & (_GEN_489 | _GEN_406);
  wire        _GEN_553 = _io_pprd_2_output != 6'h2D & (_GEN_490 | _GEN_408);
  wire        _GEN_554 = _io_pprd_2_output != 6'h2E & (_GEN_491 | _GEN_410);
  wire        _GEN_555 = _io_pprd_2_output != 6'h2F & (_GEN_492 | _GEN_412);
  wire        _GEN_556 = _io_pprd_2_output != 6'h30 & (_GEN_493 | _GEN_414);
  wire        _GEN_557 = _io_pprd_2_output != 6'h31 & (_GEN_494 | _GEN_416);
  wire        _GEN_558 = _io_pprd_2_output != 6'h32 & (_GEN_495 | _GEN_418);
  wire        _GEN_559 = _io_pprd_2_output != 6'h33 & (_GEN_496 | _GEN_420);
  wire        _GEN_560 = _io_pprd_2_output != 6'h34 & (_GEN_497 | _GEN_422);
  wire        _GEN_561 = _io_pprd_2_output != 6'h35 & (_GEN_498 | _GEN_424);
  wire        _GEN_562 = _io_pprd_2_output != 6'h36 & (_GEN_499 | _GEN_426);
  wire        _GEN_563 = _io_pprd_2_output != 6'h37 & (_GEN_500 | _GEN_428);
  wire        _GEN_564 = _io_pprd_2_output != 6'h38 & (_GEN_501 | _GEN_430);
  wire        _GEN_565 = _io_pprd_2_output != 6'h39 & (_GEN_502 | _GEN_432);
  wire        _GEN_566 = _io_pprd_2_output != 6'h3A & (_GEN_503 | _GEN_434);
  wire        _GEN_567 = _io_pprd_2_output != 6'h3B & (_GEN_504 | _GEN_436);
  wire        _GEN_568 = _io_pprd_2_output != 6'h3C & (_GEN_505 | _GEN_438);
  wire        _GEN_569 = _io_pprd_2_output != 6'h3D & (_GEN_506 | _GEN_440);
  wire        _GEN_570 = _io_pprd_2_output != 6'h3E & (_GEN_507 | _GEN_442);
  wire        _GEN_571 = _io_pprd_2_output != 6'h3F & ((&io_alloc_preg_2) | _GEN_444);
  wire        _GEN_572 = io_alloc_preg_3 == 6'h0;
  wire        _GEN_573 = io_alloc_preg_3 == 6'h1;
  wire        _GEN_574 = io_alloc_preg_3 == 6'h2;
  wire        _GEN_575 = io_alloc_preg_3 == 6'h3;
  wire        _GEN_576 = io_alloc_preg_3 == 6'h4;
  wire        _GEN_577 = io_alloc_preg_3 == 6'h5;
  wire        _GEN_578 = io_alloc_preg_3 == 6'h6;
  wire        _GEN_579 = io_alloc_preg_3 == 6'h7;
  wire        _GEN_580 = io_alloc_preg_3 == 6'h8;
  wire        _GEN_581 = io_alloc_preg_3 == 6'h9;
  wire        _GEN_582 = io_alloc_preg_3 == 6'hA;
  wire        _GEN_583 = io_alloc_preg_3 == 6'hB;
  wire        _GEN_584 = io_alloc_preg_3 == 6'hC;
  wire        _GEN_585 = io_alloc_preg_3 == 6'hD;
  wire        _GEN_586 = io_alloc_preg_3 == 6'hE;
  wire        _GEN_587 = io_alloc_preg_3 == 6'hF;
  wire        _GEN_588 = io_alloc_preg_3 == 6'h10;
  wire        _GEN_589 = io_alloc_preg_3 == 6'h11;
  wire        _GEN_590 = io_alloc_preg_3 == 6'h12;
  wire        _GEN_591 = io_alloc_preg_3 == 6'h13;
  wire        _GEN_592 = io_alloc_preg_3 == 6'h14;
  wire        _GEN_593 = io_alloc_preg_3 == 6'h15;
  wire        _GEN_594 = io_alloc_preg_3 == 6'h16;
  wire        _GEN_595 = io_alloc_preg_3 == 6'h17;
  wire        _GEN_596 = io_alloc_preg_3 == 6'h18;
  wire        _GEN_597 = io_alloc_preg_3 == 6'h19;
  wire        _GEN_598 = io_alloc_preg_3 == 6'h1A;
  wire        _GEN_599 = io_alloc_preg_3 == 6'h1B;
  wire        _GEN_600 = io_alloc_preg_3 == 6'h1C;
  wire        _GEN_601 = io_alloc_preg_3 == 6'h1D;
  wire        _GEN_602 = io_alloc_preg_3 == 6'h1E;
  wire        _GEN_603 = io_alloc_preg_3 == 6'h1F;
  wire        _GEN_604 = io_alloc_preg_3 == 6'h20;
  wire        _GEN_605 = io_alloc_preg_3 == 6'h21;
  wire        _GEN_606 = io_alloc_preg_3 == 6'h22;
  wire        _GEN_607 = io_alloc_preg_3 == 6'h23;
  wire        _GEN_608 = io_alloc_preg_3 == 6'h24;
  wire        _GEN_609 = io_alloc_preg_3 == 6'h25;
  wire        _GEN_610 = io_alloc_preg_3 == 6'h26;
  wire        _GEN_611 = io_alloc_preg_3 == 6'h27;
  wire        _GEN_612 = io_alloc_preg_3 == 6'h28;
  wire        _GEN_613 = io_alloc_preg_3 == 6'h29;
  wire        _GEN_614 = io_alloc_preg_3 == 6'h2A;
  wire        _GEN_615 = io_alloc_preg_3 == 6'h2B;
  wire        _GEN_616 = io_alloc_preg_3 == 6'h2C;
  wire        _GEN_617 = io_alloc_preg_3 == 6'h2D;
  wire        _GEN_618 = io_alloc_preg_3 == 6'h2E;
  wire        _GEN_619 = io_alloc_preg_3 == 6'h2F;
  wire        _GEN_620 = io_alloc_preg_3 == 6'h30;
  wire        _GEN_621 = io_alloc_preg_3 == 6'h31;
  wire        _GEN_622 = io_alloc_preg_3 == 6'h32;
  wire        _GEN_623 = io_alloc_preg_3 == 6'h33;
  wire        _GEN_624 = io_alloc_preg_3 == 6'h34;
  wire        _GEN_625 = io_alloc_preg_3 == 6'h35;
  wire        _GEN_626 = io_alloc_preg_3 == 6'h36;
  wire        _GEN_627 = io_alloc_preg_3 == 6'h37;
  wire        _GEN_628 = io_alloc_preg_3 == 6'h38;
  wire        _GEN_629 = io_alloc_preg_3 == 6'h39;
  wire        _GEN_630 = io_alloc_preg_3 == 6'h3A;
  wire        _GEN_631 = io_alloc_preg_3 == 6'h3B;
  wire        _GEN_632 = io_alloc_preg_3 == 6'h3C;
  wire        _GEN_633 = io_alloc_preg_3 == 6'h3D;
  wire        _GEN_634 = io_alloc_preg_3 == 6'h3E;
  always @(posedge clock) begin
    if (io_predict_fail) begin
      crat_0_valid <= io_arch_rat_0;
      crat_1_valid <= io_arch_rat_1;
      crat_2_valid <= io_arch_rat_2;
      crat_3_valid <= io_arch_rat_3;
      crat_4_valid <= io_arch_rat_4;
      crat_5_valid <= io_arch_rat_5;
      crat_6_valid <= io_arch_rat_6;
      crat_7_valid <= io_arch_rat_7;
      crat_8_valid <= io_arch_rat_8;
      crat_9_valid <= io_arch_rat_9;
      crat_10_valid <= io_arch_rat_10;
      crat_11_valid <= io_arch_rat_11;
      crat_12_valid <= io_arch_rat_12;
      crat_13_valid <= io_arch_rat_13;
      crat_14_valid <= io_arch_rat_14;
      crat_15_valid <= io_arch_rat_15;
      crat_16_valid <= io_arch_rat_16;
      crat_17_valid <= io_arch_rat_17;
      crat_18_valid <= io_arch_rat_18;
      crat_19_valid <= io_arch_rat_19;
      crat_20_valid <= io_arch_rat_20;
      crat_21_valid <= io_arch_rat_21;
      crat_22_valid <= io_arch_rat_22;
      crat_23_valid <= io_arch_rat_23;
      crat_24_valid <= io_arch_rat_24;
      crat_25_valid <= io_arch_rat_25;
      crat_26_valid <= io_arch_rat_26;
      crat_27_valid <= io_arch_rat_27;
      crat_28_valid <= io_arch_rat_28;
      crat_29_valid <= io_arch_rat_29;
      crat_30_valid <= io_arch_rat_30;
      crat_31_valid <= io_arch_rat_31;
      crat_32_valid <= io_arch_rat_32;
      crat_33_valid <= io_arch_rat_33;
      crat_34_valid <= io_arch_rat_34;
      crat_35_valid <= io_arch_rat_35;
      crat_36_valid <= io_arch_rat_36;
      crat_37_valid <= io_arch_rat_37;
      crat_38_valid <= io_arch_rat_38;
      crat_39_valid <= io_arch_rat_39;
      crat_40_valid <= io_arch_rat_40;
      crat_41_valid <= io_arch_rat_41;
      crat_42_valid <= io_arch_rat_42;
      crat_43_valid <= io_arch_rat_43;
      crat_44_valid <= io_arch_rat_44;
      crat_45_valid <= io_arch_rat_45;
      crat_46_valid <= io_arch_rat_46;
      crat_47_valid <= io_arch_rat_47;
      crat_48_valid <= io_arch_rat_48;
      crat_49_valid <= io_arch_rat_49;
      crat_50_valid <= io_arch_rat_50;
      crat_51_valid <= io_arch_rat_51;
      crat_52_valid <= io_arch_rat_52;
      crat_53_valid <= io_arch_rat_53;
      crat_54_valid <= io_arch_rat_54;
      crat_55_valid <= io_arch_rat_55;
      crat_56_valid <= io_arch_rat_56;
      crat_57_valid <= io_arch_rat_57;
      crat_58_valid <= io_arch_rat_58;
      crat_59_valid <= io_arch_rat_59;
      crat_60_valid <= io_arch_rat_60;
      crat_61_valid <= io_arch_rat_61;
      crat_62_valid <= io_arch_rat_62;
      crat_63_valid <= io_arch_rat_63;
    end
    else begin
      if (io_rd_valid_3) begin
        crat_0_valid <=
          (|_io_pprd_3_output) & (_GEN_572 | (io_rd_valid_2 ? _GEN_508 : _GEN_318));
        crat_1_valid <=
          _io_pprd_3_output != 6'h1 & (_GEN_573 | (io_rd_valid_2 ? _GEN_509 : _GEN_320));
        crat_2_valid <=
          _io_pprd_3_output != 6'h2 & (_GEN_574 | (io_rd_valid_2 ? _GEN_510 : _GEN_322));
        crat_3_valid <=
          _io_pprd_3_output != 6'h3 & (_GEN_575 | (io_rd_valid_2 ? _GEN_511 : _GEN_324));
        crat_4_valid <=
          _io_pprd_3_output != 6'h4 & (_GEN_576 | (io_rd_valid_2 ? _GEN_512 : _GEN_326));
        crat_5_valid <=
          _io_pprd_3_output != 6'h5 & (_GEN_577 | (io_rd_valid_2 ? _GEN_513 : _GEN_328));
        crat_6_valid <=
          _io_pprd_3_output != 6'h6 & (_GEN_578 | (io_rd_valid_2 ? _GEN_514 : _GEN_330));
        crat_7_valid <=
          _io_pprd_3_output != 6'h7 & (_GEN_579 | (io_rd_valid_2 ? _GEN_515 : _GEN_332));
        crat_8_valid <=
          _io_pprd_3_output != 6'h8 & (_GEN_580 | (io_rd_valid_2 ? _GEN_516 : _GEN_334));
        crat_9_valid <=
          _io_pprd_3_output != 6'h9 & (_GEN_581 | (io_rd_valid_2 ? _GEN_517 : _GEN_336));
        crat_10_valid <=
          _io_pprd_3_output != 6'hA & (_GEN_582 | (io_rd_valid_2 ? _GEN_518 : _GEN_338));
        crat_11_valid <=
          _io_pprd_3_output != 6'hB & (_GEN_583 | (io_rd_valid_2 ? _GEN_519 : _GEN_340));
        crat_12_valid <=
          _io_pprd_3_output != 6'hC & (_GEN_584 | (io_rd_valid_2 ? _GEN_520 : _GEN_342));
        crat_13_valid <=
          _io_pprd_3_output != 6'hD & (_GEN_585 | (io_rd_valid_2 ? _GEN_521 : _GEN_344));
        crat_14_valid <=
          _io_pprd_3_output != 6'hE & (_GEN_586 | (io_rd_valid_2 ? _GEN_522 : _GEN_346));
        crat_15_valid <=
          _io_pprd_3_output != 6'hF & (_GEN_587 | (io_rd_valid_2 ? _GEN_523 : _GEN_348));
        crat_16_valid <=
          _io_pprd_3_output != 6'h10 & (_GEN_588 | (io_rd_valid_2 ? _GEN_524 : _GEN_350));
        crat_17_valid <=
          _io_pprd_3_output != 6'h11 & (_GEN_589 | (io_rd_valid_2 ? _GEN_525 : _GEN_352));
        crat_18_valid <=
          _io_pprd_3_output != 6'h12 & (_GEN_590 | (io_rd_valid_2 ? _GEN_526 : _GEN_354));
        crat_19_valid <=
          _io_pprd_3_output != 6'h13 & (_GEN_591 | (io_rd_valid_2 ? _GEN_527 : _GEN_356));
        crat_20_valid <=
          _io_pprd_3_output != 6'h14 & (_GEN_592 | (io_rd_valid_2 ? _GEN_528 : _GEN_358));
        crat_21_valid <=
          _io_pprd_3_output != 6'h15 & (_GEN_593 | (io_rd_valid_2 ? _GEN_529 : _GEN_360));
        crat_22_valid <=
          _io_pprd_3_output != 6'h16 & (_GEN_594 | (io_rd_valid_2 ? _GEN_530 : _GEN_362));
        crat_23_valid <=
          _io_pprd_3_output != 6'h17 & (_GEN_595 | (io_rd_valid_2 ? _GEN_531 : _GEN_364));
        crat_24_valid <=
          _io_pprd_3_output != 6'h18 & (_GEN_596 | (io_rd_valid_2 ? _GEN_532 : _GEN_366));
        crat_25_valid <=
          _io_pprd_3_output != 6'h19 & (_GEN_597 | (io_rd_valid_2 ? _GEN_533 : _GEN_368));
        crat_26_valid <=
          _io_pprd_3_output != 6'h1A & (_GEN_598 | (io_rd_valid_2 ? _GEN_534 : _GEN_370));
        crat_27_valid <=
          _io_pprd_3_output != 6'h1B & (_GEN_599 | (io_rd_valid_2 ? _GEN_535 : _GEN_372));
        crat_28_valid <=
          _io_pprd_3_output != 6'h1C & (_GEN_600 | (io_rd_valid_2 ? _GEN_536 : _GEN_374));
        crat_29_valid <=
          _io_pprd_3_output != 6'h1D & (_GEN_601 | (io_rd_valid_2 ? _GEN_537 : _GEN_376));
        crat_30_valid <=
          _io_pprd_3_output != 6'h1E & (_GEN_602 | (io_rd_valid_2 ? _GEN_538 : _GEN_378));
        crat_31_valid <=
          _io_pprd_3_output != 6'h1F & (_GEN_603 | (io_rd_valid_2 ? _GEN_539 : _GEN_380));
        crat_32_valid <=
          _io_pprd_3_output != 6'h20 & (_GEN_604 | (io_rd_valid_2 ? _GEN_540 : _GEN_382));
        crat_33_valid <=
          _io_pprd_3_output != 6'h21 & (_GEN_605 | (io_rd_valid_2 ? _GEN_541 : _GEN_384));
        crat_34_valid <=
          _io_pprd_3_output != 6'h22 & (_GEN_606 | (io_rd_valid_2 ? _GEN_542 : _GEN_386));
        crat_35_valid <=
          _io_pprd_3_output != 6'h23 & (_GEN_607 | (io_rd_valid_2 ? _GEN_543 : _GEN_388));
        crat_36_valid <=
          _io_pprd_3_output != 6'h24 & (_GEN_608 | (io_rd_valid_2 ? _GEN_544 : _GEN_390));
        crat_37_valid <=
          _io_pprd_3_output != 6'h25 & (_GEN_609 | (io_rd_valid_2 ? _GEN_545 : _GEN_392));
        crat_38_valid <=
          _io_pprd_3_output != 6'h26 & (_GEN_610 | (io_rd_valid_2 ? _GEN_546 : _GEN_394));
        crat_39_valid <=
          _io_pprd_3_output != 6'h27 & (_GEN_611 | (io_rd_valid_2 ? _GEN_547 : _GEN_396));
        crat_40_valid <=
          _io_pprd_3_output != 6'h28 & (_GEN_612 | (io_rd_valid_2 ? _GEN_548 : _GEN_398));
        crat_41_valid <=
          _io_pprd_3_output != 6'h29 & (_GEN_613 | (io_rd_valid_2 ? _GEN_549 : _GEN_400));
        crat_42_valid <=
          _io_pprd_3_output != 6'h2A & (_GEN_614 | (io_rd_valid_2 ? _GEN_550 : _GEN_402));
        crat_43_valid <=
          _io_pprd_3_output != 6'h2B & (_GEN_615 | (io_rd_valid_2 ? _GEN_551 : _GEN_404));
        crat_44_valid <=
          _io_pprd_3_output != 6'h2C & (_GEN_616 | (io_rd_valid_2 ? _GEN_552 : _GEN_406));
        crat_45_valid <=
          _io_pprd_3_output != 6'h2D & (_GEN_617 | (io_rd_valid_2 ? _GEN_553 : _GEN_408));
        crat_46_valid <=
          _io_pprd_3_output != 6'h2E & (_GEN_618 | (io_rd_valid_2 ? _GEN_554 : _GEN_410));
        crat_47_valid <=
          _io_pprd_3_output != 6'h2F & (_GEN_619 | (io_rd_valid_2 ? _GEN_555 : _GEN_412));
        crat_48_valid <=
          _io_pprd_3_output != 6'h30 & (_GEN_620 | (io_rd_valid_2 ? _GEN_556 : _GEN_414));
        crat_49_valid <=
          _io_pprd_3_output != 6'h31 & (_GEN_621 | (io_rd_valid_2 ? _GEN_557 : _GEN_416));
        crat_50_valid <=
          _io_pprd_3_output != 6'h32 & (_GEN_622 | (io_rd_valid_2 ? _GEN_558 : _GEN_418));
        crat_51_valid <=
          _io_pprd_3_output != 6'h33 & (_GEN_623 | (io_rd_valid_2 ? _GEN_559 : _GEN_420));
        crat_52_valid <=
          _io_pprd_3_output != 6'h34 & (_GEN_624 | (io_rd_valid_2 ? _GEN_560 : _GEN_422));
        crat_53_valid <=
          _io_pprd_3_output != 6'h35 & (_GEN_625 | (io_rd_valid_2 ? _GEN_561 : _GEN_424));
        crat_54_valid <=
          _io_pprd_3_output != 6'h36 & (_GEN_626 | (io_rd_valid_2 ? _GEN_562 : _GEN_426));
        crat_55_valid <=
          _io_pprd_3_output != 6'h37 & (_GEN_627 | (io_rd_valid_2 ? _GEN_563 : _GEN_428));
        crat_56_valid <=
          _io_pprd_3_output != 6'h38 & (_GEN_628 | (io_rd_valid_2 ? _GEN_564 : _GEN_430));
        crat_57_valid <=
          _io_pprd_3_output != 6'h39 & (_GEN_629 | (io_rd_valid_2 ? _GEN_565 : _GEN_432));
        crat_58_valid <=
          _io_pprd_3_output != 6'h3A & (_GEN_630 | (io_rd_valid_2 ? _GEN_566 : _GEN_434));
        crat_59_valid <=
          _io_pprd_3_output != 6'h3B & (_GEN_631 | (io_rd_valid_2 ? _GEN_567 : _GEN_436));
        crat_60_valid <=
          _io_pprd_3_output != 6'h3C & (_GEN_632 | (io_rd_valid_2 ? _GEN_568 : _GEN_438));
        crat_61_valid <=
          _io_pprd_3_output != 6'h3D & (_GEN_633 | (io_rd_valid_2 ? _GEN_569 : _GEN_440));
        crat_62_valid <=
          _io_pprd_3_output != 6'h3E & (_GEN_634 | (io_rd_valid_2 ? _GEN_570 : _GEN_442));
        crat_63_valid <=
          _io_pprd_3_output != 6'h3F
          & ((&io_alloc_preg_3) | (io_rd_valid_2 ? _GEN_571 : _GEN_444));
      end
      else if (io_rd_valid_2) begin
        crat_0_valid <= _GEN_508;
        crat_1_valid <= _GEN_509;
        crat_2_valid <= _GEN_510;
        crat_3_valid <= _GEN_511;
        crat_4_valid <= _GEN_512;
        crat_5_valid <= _GEN_513;
        crat_6_valid <= _GEN_514;
        crat_7_valid <= _GEN_515;
        crat_8_valid <= _GEN_516;
        crat_9_valid <= _GEN_517;
        crat_10_valid <= _GEN_518;
        crat_11_valid <= _GEN_519;
        crat_12_valid <= _GEN_520;
        crat_13_valid <= _GEN_521;
        crat_14_valid <= _GEN_522;
        crat_15_valid <= _GEN_523;
        crat_16_valid <= _GEN_524;
        crat_17_valid <= _GEN_525;
        crat_18_valid <= _GEN_526;
        crat_19_valid <= _GEN_527;
        crat_20_valid <= _GEN_528;
        crat_21_valid <= _GEN_529;
        crat_22_valid <= _GEN_530;
        crat_23_valid <= _GEN_531;
        crat_24_valid <= _GEN_532;
        crat_25_valid <= _GEN_533;
        crat_26_valid <= _GEN_534;
        crat_27_valid <= _GEN_535;
        crat_28_valid <= _GEN_536;
        crat_29_valid <= _GEN_537;
        crat_30_valid <= _GEN_538;
        crat_31_valid <= _GEN_539;
        crat_32_valid <= _GEN_540;
        crat_33_valid <= _GEN_541;
        crat_34_valid <= _GEN_542;
        crat_35_valid <= _GEN_543;
        crat_36_valid <= _GEN_544;
        crat_37_valid <= _GEN_545;
        crat_38_valid <= _GEN_546;
        crat_39_valid <= _GEN_547;
        crat_40_valid <= _GEN_548;
        crat_41_valid <= _GEN_549;
        crat_42_valid <= _GEN_550;
        crat_43_valid <= _GEN_551;
        crat_44_valid <= _GEN_552;
        crat_45_valid <= _GEN_553;
        crat_46_valid <= _GEN_554;
        crat_47_valid <= _GEN_555;
        crat_48_valid <= _GEN_556;
        crat_49_valid <= _GEN_557;
        crat_50_valid <= _GEN_558;
        crat_51_valid <= _GEN_559;
        crat_52_valid <= _GEN_560;
        crat_53_valid <= _GEN_561;
        crat_54_valid <= _GEN_562;
        crat_55_valid <= _GEN_563;
        crat_56_valid <= _GEN_564;
        crat_57_valid <= _GEN_565;
        crat_58_valid <= _GEN_566;
        crat_59_valid <= _GEN_567;
        crat_60_valid <= _GEN_568;
        crat_61_valid <= _GEN_569;
        crat_62_valid <= _GEN_570;
        crat_63_valid <= _GEN_571;
      end
      else if (io_rd_valid_1) begin
        crat_0_valid <= _GEN_317;
        crat_1_valid <= _GEN_319;
        crat_2_valid <= _GEN_321;
        crat_3_valid <= _GEN_323;
        crat_4_valid <= _GEN_325;
        crat_5_valid <= _GEN_327;
        crat_6_valid <= _GEN_329;
        crat_7_valid <= _GEN_331;
        crat_8_valid <= _GEN_333;
        crat_9_valid <= _GEN_335;
        crat_10_valid <= _GEN_337;
        crat_11_valid <= _GEN_339;
        crat_12_valid <= _GEN_341;
        crat_13_valid <= _GEN_343;
        crat_14_valid <= _GEN_345;
        crat_15_valid <= _GEN_347;
        crat_16_valid <= _GEN_349;
        crat_17_valid <= _GEN_351;
        crat_18_valid <= _GEN_353;
        crat_19_valid <= _GEN_355;
        crat_20_valid <= _GEN_357;
        crat_21_valid <= _GEN_359;
        crat_22_valid <= _GEN_361;
        crat_23_valid <= _GEN_363;
        crat_24_valid <= _GEN_365;
        crat_25_valid <= _GEN_367;
        crat_26_valid <= _GEN_369;
        crat_27_valid <= _GEN_371;
        crat_28_valid <= _GEN_373;
        crat_29_valid <= _GEN_375;
        crat_30_valid <= _GEN_377;
        crat_31_valid <= _GEN_379;
        crat_32_valid <= _GEN_381;
        crat_33_valid <= _GEN_383;
        crat_34_valid <= _GEN_385;
        crat_35_valid <= _GEN_387;
        crat_36_valid <= _GEN_389;
        crat_37_valid <= _GEN_391;
        crat_38_valid <= _GEN_393;
        crat_39_valid <= _GEN_395;
        crat_40_valid <= _GEN_397;
        crat_41_valid <= _GEN_399;
        crat_42_valid <= _GEN_401;
        crat_43_valid <= _GEN_403;
        crat_44_valid <= _GEN_405;
        crat_45_valid <= _GEN_407;
        crat_46_valid <= _GEN_409;
        crat_47_valid <= _GEN_411;
        crat_48_valid <= _GEN_413;
        crat_49_valid <= _GEN_415;
        crat_50_valid <= _GEN_417;
        crat_51_valid <= _GEN_419;
        crat_52_valid <= _GEN_421;
        crat_53_valid <= _GEN_423;
        crat_54_valid <= _GEN_425;
        crat_55_valid <= _GEN_427;
        crat_56_valid <= _GEN_429;
        crat_57_valid <= _GEN_431;
        crat_58_valid <= _GEN_433;
        crat_59_valid <= _GEN_435;
        crat_60_valid <= _GEN_437;
        crat_61_valid <= _GEN_439;
        crat_62_valid <= _GEN_441;
        crat_63_valid <= _GEN_443;
      end
      else if (io_rd_valid_0) begin
        crat_0_valid <= _GEN_126;
        crat_1_valid <= _GEN_128;
        crat_2_valid <= _GEN_130;
        crat_3_valid <= _GEN_132;
        crat_4_valid <= _GEN_134;
        crat_5_valid <= _GEN_136;
        crat_6_valid <= _GEN_138;
        crat_7_valid <= _GEN_140;
        crat_8_valid <= _GEN_142;
        crat_9_valid <= _GEN_144;
        crat_10_valid <= _GEN_146;
        crat_11_valid <= _GEN_148;
        crat_12_valid <= _GEN_150;
        crat_13_valid <= _GEN_152;
        crat_14_valid <= _GEN_154;
        crat_15_valid <= _GEN_156;
        crat_16_valid <= _GEN_158;
        crat_17_valid <= _GEN_160;
        crat_18_valid <= _GEN_162;
        crat_19_valid <= _GEN_164;
        crat_20_valid <= _GEN_166;
        crat_21_valid <= _GEN_168;
        crat_22_valid <= _GEN_170;
        crat_23_valid <= _GEN_172;
        crat_24_valid <= _GEN_174;
        crat_25_valid <= _GEN_176;
        crat_26_valid <= _GEN_178;
        crat_27_valid <= _GEN_180;
        crat_28_valid <= _GEN_182;
        crat_29_valid <= _GEN_184;
        crat_30_valid <= _GEN_186;
        crat_31_valid <= _GEN_188;
        crat_32_valid <= _GEN_190;
        crat_33_valid <= _GEN_192;
        crat_34_valid <= _GEN_194;
        crat_35_valid <= _GEN_196;
        crat_36_valid <= _GEN_198;
        crat_37_valid <= _GEN_200;
        crat_38_valid <= _GEN_202;
        crat_39_valid <= _GEN_204;
        crat_40_valid <= _GEN_206;
        crat_41_valid <= _GEN_208;
        crat_42_valid <= _GEN_210;
        crat_43_valid <= _GEN_212;
        crat_44_valid <= _GEN_214;
        crat_45_valid <= _GEN_216;
        crat_46_valid <= _GEN_218;
        crat_47_valid <= _GEN_220;
        crat_48_valid <= _GEN_222;
        crat_49_valid <= _GEN_224;
        crat_50_valid <= _GEN_226;
        crat_51_valid <= _GEN_228;
        crat_52_valid <= _GEN_230;
        crat_53_valid <= _GEN_232;
        crat_54_valid <= _GEN_234;
        crat_55_valid <= _GEN_236;
        crat_56_valid <= _GEN_238;
        crat_57_valid <= _GEN_240;
        crat_58_valid <= _GEN_242;
        crat_59_valid <= _GEN_244;
        crat_60_valid <= _GEN_246;
        crat_61_valid <= _GEN_248;
        crat_62_valid <= _GEN_250;
        crat_63_valid <= _GEN_252;
      end
      else begin
        crat_0_valid <= _GEN;
        crat_1_valid <= _GEN_0;
        crat_2_valid <= _GEN_1;
        crat_3_valid <= _GEN_2;
        crat_4_valid <= _GEN_3;
        crat_5_valid <= _GEN_4;
        crat_6_valid <= _GEN_5;
        crat_7_valid <= _GEN_6;
        crat_8_valid <= _GEN_7;
        crat_9_valid <= _GEN_8;
        crat_10_valid <= _GEN_9;
        crat_11_valid <= _GEN_10;
        crat_12_valid <= _GEN_11;
        crat_13_valid <= _GEN_12;
        crat_14_valid <= _GEN_13;
        crat_15_valid <= _GEN_14;
        crat_16_valid <= _GEN_15;
        crat_17_valid <= _GEN_16;
        crat_18_valid <= _GEN_17;
        crat_19_valid <= _GEN_18;
        crat_20_valid <= _GEN_19;
        crat_21_valid <= _GEN_20;
        crat_22_valid <= _GEN_21;
        crat_23_valid <= _GEN_22;
        crat_24_valid <= _GEN_23;
        crat_25_valid <= _GEN_24;
        crat_26_valid <= _GEN_25;
        crat_27_valid <= _GEN_26;
        crat_28_valid <= _GEN_27;
        crat_29_valid <= _GEN_28;
        crat_30_valid <= _GEN_29;
        crat_31_valid <= _GEN_30;
        crat_32_valid <= _GEN_31;
        crat_33_valid <= _GEN_32;
        crat_34_valid <= _GEN_33;
        crat_35_valid <= _GEN_34;
        crat_36_valid <= _GEN_35;
        crat_37_valid <= _GEN_36;
        crat_38_valid <= _GEN_37;
        crat_39_valid <= _GEN_38;
        crat_40_valid <= _GEN_39;
        crat_41_valid <= _GEN_40;
        crat_42_valid <= _GEN_41;
        crat_43_valid <= _GEN_42;
        crat_44_valid <= _GEN_43;
        crat_45_valid <= _GEN_44;
        crat_46_valid <= _GEN_45;
        crat_47_valid <= _GEN_46;
        crat_48_valid <= _GEN_47;
        crat_49_valid <= _GEN_48;
        crat_50_valid <= _GEN_49;
        crat_51_valid <= _GEN_50;
        crat_52_valid <= _GEN_51;
        crat_53_valid <= _GEN_52;
        crat_54_valid <= _GEN_53;
        crat_55_valid <= _GEN_54;
        crat_56_valid <= _GEN_55;
        crat_57_valid <= _GEN_56;
        crat_58_valid <= _GEN_57;
        crat_59_valid <= _GEN_58;
        crat_60_valid <= _GEN_59;
        crat_61_valid <= _GEN_60;
        crat_62_valid <= _GEN_61;
        crat_63_valid <= _GEN_62;
      end
      if (io_rd_valid_3 & _GEN_572)
        crat_0_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_445)
        crat_0_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_254)
        crat_0_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_63)
        crat_0_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_573)
        crat_1_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_446)
        crat_1_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_255)
        crat_1_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_64)
        crat_1_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_574)
        crat_2_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_447)
        crat_2_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_256)
        crat_2_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_65)
        crat_2_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_575)
        crat_3_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_448)
        crat_3_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_257)
        crat_3_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_66)
        crat_3_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_576)
        crat_4_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_449)
        crat_4_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_258)
        crat_4_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_67)
        crat_4_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_577)
        crat_5_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_450)
        crat_5_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_259)
        crat_5_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_68)
        crat_5_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_578)
        crat_6_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_451)
        crat_6_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_260)
        crat_6_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_69)
        crat_6_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_579)
        crat_7_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_452)
        crat_7_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_261)
        crat_7_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_70)
        crat_7_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_580)
        crat_8_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_453)
        crat_8_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_262)
        crat_8_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_71)
        crat_8_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_581)
        crat_9_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_454)
        crat_9_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_263)
        crat_9_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_72)
        crat_9_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_582)
        crat_10_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_455)
        crat_10_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_264)
        crat_10_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_73)
        crat_10_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_583)
        crat_11_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_456)
        crat_11_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_265)
        crat_11_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_74)
        crat_11_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_584)
        crat_12_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_457)
        crat_12_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_266)
        crat_12_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_75)
        crat_12_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_585)
        crat_13_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_458)
        crat_13_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_267)
        crat_13_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_76)
        crat_13_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_586)
        crat_14_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_459)
        crat_14_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_268)
        crat_14_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_77)
        crat_14_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_587)
        crat_15_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_460)
        crat_15_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_269)
        crat_15_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_78)
        crat_15_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_588)
        crat_16_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_461)
        crat_16_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_270)
        crat_16_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_79)
        crat_16_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_589)
        crat_17_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_462)
        crat_17_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_271)
        crat_17_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_80)
        crat_17_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_590)
        crat_18_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_463)
        crat_18_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_272)
        crat_18_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_81)
        crat_18_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_591)
        crat_19_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_464)
        crat_19_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_273)
        crat_19_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_82)
        crat_19_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_592)
        crat_20_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_465)
        crat_20_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_274)
        crat_20_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_83)
        crat_20_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_593)
        crat_21_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_466)
        crat_21_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_275)
        crat_21_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_84)
        crat_21_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_594)
        crat_22_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_467)
        crat_22_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_276)
        crat_22_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_85)
        crat_22_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_595)
        crat_23_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_468)
        crat_23_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_277)
        crat_23_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_86)
        crat_23_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_596)
        crat_24_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_469)
        crat_24_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_278)
        crat_24_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_87)
        crat_24_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_597)
        crat_25_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_470)
        crat_25_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_279)
        crat_25_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_88)
        crat_25_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_598)
        crat_26_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_471)
        crat_26_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_280)
        crat_26_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_89)
        crat_26_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_599)
        crat_27_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_472)
        crat_27_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_281)
        crat_27_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_90)
        crat_27_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_600)
        crat_28_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_473)
        crat_28_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_282)
        crat_28_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_91)
        crat_28_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_601)
        crat_29_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_474)
        crat_29_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_283)
        crat_29_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_92)
        crat_29_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_602)
        crat_30_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_475)
        crat_30_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_284)
        crat_30_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_93)
        crat_30_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_603)
        crat_31_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_476)
        crat_31_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_285)
        crat_31_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_94)
        crat_31_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_604)
        crat_32_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_477)
        crat_32_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_286)
        crat_32_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_95)
        crat_32_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_605)
        crat_33_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_478)
        crat_33_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_287)
        crat_33_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_96)
        crat_33_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_606)
        crat_34_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_479)
        crat_34_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_288)
        crat_34_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_97)
        crat_34_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_607)
        crat_35_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_480)
        crat_35_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_289)
        crat_35_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_98)
        crat_35_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_608)
        crat_36_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_481)
        crat_36_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_290)
        crat_36_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_99)
        crat_36_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_609)
        crat_37_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_482)
        crat_37_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_291)
        crat_37_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_100)
        crat_37_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_610)
        crat_38_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_483)
        crat_38_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_292)
        crat_38_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_101)
        crat_38_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_611)
        crat_39_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_484)
        crat_39_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_293)
        crat_39_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_102)
        crat_39_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_612)
        crat_40_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_485)
        crat_40_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_294)
        crat_40_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_103)
        crat_40_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_613)
        crat_41_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_486)
        crat_41_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_295)
        crat_41_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_104)
        crat_41_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_614)
        crat_42_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_487)
        crat_42_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_296)
        crat_42_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_105)
        crat_42_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_615)
        crat_43_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_488)
        crat_43_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_297)
        crat_43_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_106)
        crat_43_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_616)
        crat_44_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_489)
        crat_44_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_298)
        crat_44_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_107)
        crat_44_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_617)
        crat_45_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_490)
        crat_45_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_299)
        crat_45_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_108)
        crat_45_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_618)
        crat_46_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_491)
        crat_46_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_300)
        crat_46_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_109)
        crat_46_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_619)
        crat_47_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_492)
        crat_47_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_301)
        crat_47_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_110)
        crat_47_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_620)
        crat_48_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_493)
        crat_48_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_302)
        crat_48_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_111)
        crat_48_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_621)
        crat_49_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_494)
        crat_49_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_303)
        crat_49_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_112)
        crat_49_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_622)
        crat_50_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_495)
        crat_50_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_304)
        crat_50_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_113)
        crat_50_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_623)
        crat_51_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_496)
        crat_51_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_305)
        crat_51_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_114)
        crat_51_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_624)
        crat_52_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_497)
        crat_52_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_306)
        crat_52_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_115)
        crat_52_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_625)
        crat_53_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_498)
        crat_53_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_307)
        crat_53_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_116)
        crat_53_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_626)
        crat_54_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_499)
        crat_54_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_308)
        crat_54_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_117)
        crat_54_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_627)
        crat_55_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_500)
        crat_55_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_309)
        crat_55_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_118)
        crat_55_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_628)
        crat_56_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_501)
        crat_56_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_310)
        crat_56_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_119)
        crat_56_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_629)
        crat_57_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_502)
        crat_57_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_311)
        crat_57_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_120)
        crat_57_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_630)
        crat_58_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_503)
        crat_58_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_312)
        crat_58_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_121)
        crat_58_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_631)
        crat_59_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_504)
        crat_59_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_313)
        crat_59_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_122)
        crat_59_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_632)
        crat_60_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_505)
        crat_60_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_314)
        crat_60_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_123)
        crat_60_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_633)
        crat_61_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_506)
        crat_61_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_315)
        crat_61_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_124)
        crat_61_lr <= io_rd_0;
      if (io_rd_valid_3 & _GEN_634)
        crat_62_lr <= io_rd_3;
      else if (io_rd_valid_2 & _GEN_507)
        crat_62_lr <= io_rd_2;
      else if (io_rd_valid_1 & _GEN_316)
        crat_62_lr <= io_rd_1;
      else if (io_rd_valid_0 & _GEN_125)
        crat_62_lr <= io_rd_0;
      if (io_rd_valid_3 & (&io_alloc_preg_3))
        crat_63_lr <= io_rd_3;
      else if (io_rd_valid_2 & (&io_alloc_preg_2))
        crat_63_lr <= io_rd_2;
      else if (io_rd_valid_1 & (&io_alloc_preg_1))
        crat_63_lr <= io_rd_1;
      else if (io_rd_valid_0 & (&io_alloc_preg_0))
        crat_63_lr <= io_rd_0;
    end
  end // always @(posedge)
  assign io_prj_0 =
    {|{rj_hit_oh_0_63,
       rj_hit_oh_0_62,
       rj_hit_oh_0_61,
       rj_hit_oh_0_60,
       rj_hit_oh_0_59,
       rj_hit_oh_0_58,
       rj_hit_oh_0_57,
       rj_hit_oh_0_56,
       rj_hit_oh_0_55,
       rj_hit_oh_0_54,
       rj_hit_oh_0_53,
       rj_hit_oh_0_52,
       rj_hit_oh_0_51,
       rj_hit_oh_0_50,
       rj_hit_oh_0_49,
       rj_hit_oh_0_48,
       rj_hit_oh_0_47,
       rj_hit_oh_0_46,
       rj_hit_oh_0_45,
       rj_hit_oh_0_44,
       rj_hit_oh_0_43,
       rj_hit_oh_0_42,
       rj_hit_oh_0_41,
       rj_hit_oh_0_40,
       rj_hit_oh_0_39,
       rj_hit_oh_0_38,
       rj_hit_oh_0_37,
       rj_hit_oh_0_36,
       rj_hit_oh_0_35,
       rj_hit_oh_0_34,
       rj_hit_oh_0_33,
       crat_32_valid & crat_32_lr == io_rj_0},
     |(_io_prj_0_T_1073[30:15]),
     |(_io_prj_0_T_1075[14:7]),
     |(_io_prj_0_T_1077[6:3]),
     |(_io_prj_0_T_1079[2:1]),
     _io_prj_0_T_1079[2] | _io_prj_0_T_1079[0]};
  assign io_prj_1 =
    {|{rj_hit_oh_1_63,
       rj_hit_oh_1_62,
       rj_hit_oh_1_61,
       rj_hit_oh_1_60,
       rj_hit_oh_1_59,
       rj_hit_oh_1_58,
       rj_hit_oh_1_57,
       rj_hit_oh_1_56,
       rj_hit_oh_1_55,
       rj_hit_oh_1_54,
       rj_hit_oh_1_53,
       rj_hit_oh_1_52,
       rj_hit_oh_1_51,
       rj_hit_oh_1_50,
       rj_hit_oh_1_49,
       rj_hit_oh_1_48,
       rj_hit_oh_1_47,
       rj_hit_oh_1_46,
       rj_hit_oh_1_45,
       rj_hit_oh_1_44,
       rj_hit_oh_1_43,
       rj_hit_oh_1_42,
       rj_hit_oh_1_41,
       rj_hit_oh_1_40,
       rj_hit_oh_1_39,
       rj_hit_oh_1_38,
       rj_hit_oh_1_37,
       rj_hit_oh_1_36,
       rj_hit_oh_1_35,
       rj_hit_oh_1_34,
       rj_hit_oh_1_33,
       crat_32_valid & crat_32_lr == io_rj_1},
     |(_io_prj_1_T_1073[30:15]),
     |(_io_prj_1_T_1075[14:7]),
     |(_io_prj_1_T_1077[6:3]),
     |(_io_prj_1_T_1079[2:1]),
     _io_prj_1_T_1079[2] | _io_prj_1_T_1079[0]};
  assign io_prj_2 =
    {|{rj_hit_oh_2_63,
       rj_hit_oh_2_62,
       rj_hit_oh_2_61,
       rj_hit_oh_2_60,
       rj_hit_oh_2_59,
       rj_hit_oh_2_58,
       rj_hit_oh_2_57,
       rj_hit_oh_2_56,
       rj_hit_oh_2_55,
       rj_hit_oh_2_54,
       rj_hit_oh_2_53,
       rj_hit_oh_2_52,
       rj_hit_oh_2_51,
       rj_hit_oh_2_50,
       rj_hit_oh_2_49,
       rj_hit_oh_2_48,
       rj_hit_oh_2_47,
       rj_hit_oh_2_46,
       rj_hit_oh_2_45,
       rj_hit_oh_2_44,
       rj_hit_oh_2_43,
       rj_hit_oh_2_42,
       rj_hit_oh_2_41,
       rj_hit_oh_2_40,
       rj_hit_oh_2_39,
       rj_hit_oh_2_38,
       rj_hit_oh_2_37,
       rj_hit_oh_2_36,
       rj_hit_oh_2_35,
       rj_hit_oh_2_34,
       rj_hit_oh_2_33,
       crat_32_valid & crat_32_lr == io_rj_2},
     |(_io_prj_2_T_1073[30:15]),
     |(_io_prj_2_T_1075[14:7]),
     |(_io_prj_2_T_1077[6:3]),
     |(_io_prj_2_T_1079[2:1]),
     _io_prj_2_T_1079[2] | _io_prj_2_T_1079[0]};
  assign io_prj_3 =
    {|{rj_hit_oh_3_63,
       rj_hit_oh_3_62,
       rj_hit_oh_3_61,
       rj_hit_oh_3_60,
       rj_hit_oh_3_59,
       rj_hit_oh_3_58,
       rj_hit_oh_3_57,
       rj_hit_oh_3_56,
       rj_hit_oh_3_55,
       rj_hit_oh_3_54,
       rj_hit_oh_3_53,
       rj_hit_oh_3_52,
       rj_hit_oh_3_51,
       rj_hit_oh_3_50,
       rj_hit_oh_3_49,
       rj_hit_oh_3_48,
       rj_hit_oh_3_47,
       rj_hit_oh_3_46,
       rj_hit_oh_3_45,
       rj_hit_oh_3_44,
       rj_hit_oh_3_43,
       rj_hit_oh_3_42,
       rj_hit_oh_3_41,
       rj_hit_oh_3_40,
       rj_hit_oh_3_39,
       rj_hit_oh_3_38,
       rj_hit_oh_3_37,
       rj_hit_oh_3_36,
       rj_hit_oh_3_35,
       rj_hit_oh_3_34,
       rj_hit_oh_3_33,
       crat_32_valid & crat_32_lr == io_rj_3},
     |(_io_prj_3_T_1073[30:15]),
     |(_io_prj_3_T_1075[14:7]),
     |(_io_prj_3_T_1077[6:3]),
     |(_io_prj_3_T_1079[2:1]),
     _io_prj_3_T_1079[2] | _io_prj_3_T_1079[0]};
  assign io_prk_0 =
    {|{rk_hit_oh_0_63,
       rk_hit_oh_0_62,
       rk_hit_oh_0_61,
       rk_hit_oh_0_60,
       rk_hit_oh_0_59,
       rk_hit_oh_0_58,
       rk_hit_oh_0_57,
       rk_hit_oh_0_56,
       rk_hit_oh_0_55,
       rk_hit_oh_0_54,
       rk_hit_oh_0_53,
       rk_hit_oh_0_52,
       rk_hit_oh_0_51,
       rk_hit_oh_0_50,
       rk_hit_oh_0_49,
       rk_hit_oh_0_48,
       rk_hit_oh_0_47,
       rk_hit_oh_0_46,
       rk_hit_oh_0_45,
       rk_hit_oh_0_44,
       rk_hit_oh_0_43,
       rk_hit_oh_0_42,
       rk_hit_oh_0_41,
       rk_hit_oh_0_40,
       rk_hit_oh_0_39,
       rk_hit_oh_0_38,
       rk_hit_oh_0_37,
       rk_hit_oh_0_36,
       rk_hit_oh_0_35,
       rk_hit_oh_0_34,
       rk_hit_oh_0_33,
       crat_32_valid & crat_32_lr == io_rk_0},
     |(_io_prk_0_T_1073[30:15]),
     |(_io_prk_0_T_1075[14:7]),
     |(_io_prk_0_T_1077[6:3]),
     |(_io_prk_0_T_1079[2:1]),
     _io_prk_0_T_1079[2] | _io_prk_0_T_1079[0]};
  assign io_prk_1 =
    {|{rk_hit_oh_1_63,
       rk_hit_oh_1_62,
       rk_hit_oh_1_61,
       rk_hit_oh_1_60,
       rk_hit_oh_1_59,
       rk_hit_oh_1_58,
       rk_hit_oh_1_57,
       rk_hit_oh_1_56,
       rk_hit_oh_1_55,
       rk_hit_oh_1_54,
       rk_hit_oh_1_53,
       rk_hit_oh_1_52,
       rk_hit_oh_1_51,
       rk_hit_oh_1_50,
       rk_hit_oh_1_49,
       rk_hit_oh_1_48,
       rk_hit_oh_1_47,
       rk_hit_oh_1_46,
       rk_hit_oh_1_45,
       rk_hit_oh_1_44,
       rk_hit_oh_1_43,
       rk_hit_oh_1_42,
       rk_hit_oh_1_41,
       rk_hit_oh_1_40,
       rk_hit_oh_1_39,
       rk_hit_oh_1_38,
       rk_hit_oh_1_37,
       rk_hit_oh_1_36,
       rk_hit_oh_1_35,
       rk_hit_oh_1_34,
       rk_hit_oh_1_33,
       crat_32_valid & crat_32_lr == io_rk_1},
     |(_io_prk_1_T_1073[30:15]),
     |(_io_prk_1_T_1075[14:7]),
     |(_io_prk_1_T_1077[6:3]),
     |(_io_prk_1_T_1079[2:1]),
     _io_prk_1_T_1079[2] | _io_prk_1_T_1079[0]};
  assign io_prk_2 =
    {|{rk_hit_oh_2_63,
       rk_hit_oh_2_62,
       rk_hit_oh_2_61,
       rk_hit_oh_2_60,
       rk_hit_oh_2_59,
       rk_hit_oh_2_58,
       rk_hit_oh_2_57,
       rk_hit_oh_2_56,
       rk_hit_oh_2_55,
       rk_hit_oh_2_54,
       rk_hit_oh_2_53,
       rk_hit_oh_2_52,
       rk_hit_oh_2_51,
       rk_hit_oh_2_50,
       rk_hit_oh_2_49,
       rk_hit_oh_2_48,
       rk_hit_oh_2_47,
       rk_hit_oh_2_46,
       rk_hit_oh_2_45,
       rk_hit_oh_2_44,
       rk_hit_oh_2_43,
       rk_hit_oh_2_42,
       rk_hit_oh_2_41,
       rk_hit_oh_2_40,
       rk_hit_oh_2_39,
       rk_hit_oh_2_38,
       rk_hit_oh_2_37,
       rk_hit_oh_2_36,
       rk_hit_oh_2_35,
       rk_hit_oh_2_34,
       rk_hit_oh_2_33,
       crat_32_valid & crat_32_lr == io_rk_2},
     |(_io_prk_2_T_1073[30:15]),
     |(_io_prk_2_T_1075[14:7]),
     |(_io_prk_2_T_1077[6:3]),
     |(_io_prk_2_T_1079[2:1]),
     _io_prk_2_T_1079[2] | _io_prk_2_T_1079[0]};
  assign io_prk_3 =
    {|{rk_hit_oh_3_63,
       rk_hit_oh_3_62,
       rk_hit_oh_3_61,
       rk_hit_oh_3_60,
       rk_hit_oh_3_59,
       rk_hit_oh_3_58,
       rk_hit_oh_3_57,
       rk_hit_oh_3_56,
       rk_hit_oh_3_55,
       rk_hit_oh_3_54,
       rk_hit_oh_3_53,
       rk_hit_oh_3_52,
       rk_hit_oh_3_51,
       rk_hit_oh_3_50,
       rk_hit_oh_3_49,
       rk_hit_oh_3_48,
       rk_hit_oh_3_47,
       rk_hit_oh_3_46,
       rk_hit_oh_3_45,
       rk_hit_oh_3_44,
       rk_hit_oh_3_43,
       rk_hit_oh_3_42,
       rk_hit_oh_3_41,
       rk_hit_oh_3_40,
       rk_hit_oh_3_39,
       rk_hit_oh_3_38,
       rk_hit_oh_3_37,
       rk_hit_oh_3_36,
       rk_hit_oh_3_35,
       rk_hit_oh_3_34,
       rk_hit_oh_3_33,
       crat_32_valid & crat_32_lr == io_rk_3},
     |(_io_prk_3_T_1073[30:15]),
     |(_io_prk_3_T_1075[14:7]),
     |(_io_prk_3_T_1077[6:3]),
     |(_io_prk_3_T_1079[2:1]),
     _io_prk_3_T_1079[2] | _io_prk_3_T_1079[0]};
  assign io_pprd_0 = _io_pprd_0_output;
  assign io_pprd_1 = _io_pprd_1_output;
  assign io_pprd_2 = _io_pprd_2_output;
  assign io_pprd_3 = _io_pprd_3_output;
endmodule
